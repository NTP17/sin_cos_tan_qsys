-- megafunction wizard: %ALTFP_SINCOS%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altfp_sincos 

-- ============================================================
-- File Name: sinhw.vhd
-- Megafunction Name(s):
-- 			altfp_sincos
--
-- Simulation Library Files(s):
-- 			
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


--altfp_sincos CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" OPERATION="SIN" PIPELINE=36 ROUNDING="TO_NEAREST" WIDTH_EXP=8 WIDTH_MAN=23 clock data result
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END


--altfp_sincos_cordic_m CBX_AUTO_BLACKBOX="ALL" DEPTH=18 DEVICE_FAMILY="Cyclone V" INDEXPOINT=2 WIDTH=34 aclr clken clock indexbit radians sincos sincosbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=0 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_45b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_45b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_45b IS

	 SIGNAL  wire_cata_0_cordic_atan_w_lg_w_lg_indexbit10924w10925w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_0_cordic_atan_w_lg_indexbit10922w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_0_cordic_atan_w_lg_indexbit10924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_0_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_2_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_0_cordic_atan_w_valuenode_0_w_range10923w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_0_cordic_atan_w_valuenode_2_w_range10921w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_0_cordic_atan_w_lg_w_lg_indexbit10924w10925w(i) <= wire_cata_0_cordic_atan_w_lg_indexbit10924w(0) AND wire_cata_0_cordic_atan_w_valuenode_0_w_range10923w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_0_cordic_atan_w_lg_indexbit10922w(i) <= indexbit AND wire_cata_0_cordic_atan_w_valuenode_2_w_range10921w(i);
	END GENERATE loop1;
	wire_cata_0_cordic_atan_w_lg_indexbit10924w(0) <= NOT indexbit;
	arctan <= (wire_cata_0_cordic_atan_w_lg_w_lg_indexbit10924w10925w OR wire_cata_0_cordic_atan_w_lg_indexbit10922w);
	valuenode_0_w <= "001100100100001111110110101010001000100001011010";
	valuenode_2_w <= "000011111010110110111010111111001001011001000000";
	wire_cata_0_cordic_atan_w_valuenode_0_w_range10923w <= valuenode_0_w(47 DOWNTO 14);
	wire_cata_0_cordic_atan_w_valuenode_2_w_range10921w <= valuenode_2_w(45 DOWNTO 12);

 END RTL; --sinhw_altfp_sincos_cordic_atan_45b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=10 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_l6b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_l6b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_l6b IS

	 SIGNAL  wire_cata_10_cordic_atan_w_lg_w_lg_indexbit10930w10931w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_w_lg_indexbit10928w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_w_lg_indexbit10930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_10_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_12_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_w_valuenode_10_w_range10929w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_w_valuenode_12_w_range10927w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop2 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_10_cordic_atan_w_lg_w_lg_indexbit10930w10931w(i) <= wire_cata_10_cordic_atan_w_lg_indexbit10930w(0) AND wire_cata_10_cordic_atan_w_valuenode_10_w_range10929w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_10_cordic_atan_w_lg_indexbit10928w(i) <= indexbit AND wire_cata_10_cordic_atan_w_valuenode_12_w_range10927w(i);
	END GENERATE loop3;
	wire_cata_10_cordic_atan_w_lg_indexbit10930w(0) <= NOT indexbit;
	arctan <= (wire_cata_10_cordic_atan_w_lg_w_lg_indexbit10930w10931w OR wire_cata_10_cordic_atan_w_lg_indexbit10928w);
	valuenode_10_w <= "000000000000111111111111111111111010101010101011";
	valuenode_12_w <= "000000000000001111111111111111111111111010101011";
	wire_cata_10_cordic_atan_w_valuenode_10_w_range10929w <= valuenode_10_w(47 DOWNTO 14);
	wire_cata_10_cordic_atan_w_valuenode_12_w_range10927w <= valuenode_12_w(45 DOWNTO 12);

 END RTL; --sinhw_altfp_sincos_cordic_atan_l6b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=11 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_m6b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_m6b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_m6b IS

	 SIGNAL  wire_cata_11_cordic_atan_w_lg_w_lg_indexbit10936w10937w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_w_lg_indexbit10934w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_w_lg_indexbit10936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_11_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_13_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_w_valuenode_11_w_range10935w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_w_valuenode_13_w_range10933w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop4 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_11_cordic_atan_w_lg_w_lg_indexbit10936w10937w(i) <= wire_cata_11_cordic_atan_w_lg_indexbit10936w(0) AND wire_cata_11_cordic_atan_w_valuenode_11_w_range10935w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_11_cordic_atan_w_lg_indexbit10934w(i) <= indexbit AND wire_cata_11_cordic_atan_w_valuenode_13_w_range10933w(i);
	END GENERATE loop5;
	wire_cata_11_cordic_atan_w_lg_indexbit10936w(0) <= NOT indexbit;
	arctan <= (wire_cata_11_cordic_atan_w_lg_w_lg_indexbit10936w10937w OR wire_cata_11_cordic_atan_w_lg_indexbit10934w);
	valuenode_11_w <= "000000000000011111111111111111111111010101010101";
	valuenode_13_w <= "000000000000000111111111111111111111111111010101";
	wire_cata_11_cordic_atan_w_valuenode_11_w_range10935w <= valuenode_11_w(47 DOWNTO 14);
	wire_cata_11_cordic_atan_w_valuenode_13_w_range10933w <= valuenode_13_w(45 DOWNTO 12);

 END RTL; --sinhw_altfp_sincos_cordic_atan_m6b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=12 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_n6b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_n6b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_n6b IS

	 SIGNAL  wire_cata_12_cordic_atan_w_lg_w_lg_indexbit10942w10943w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_w_lg_indexbit10940w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_w_lg_indexbit10942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_12_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_14_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_w_valuenode_12_w_range10941w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_w_valuenode_14_w_range10939w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop6 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_12_cordic_atan_w_lg_w_lg_indexbit10942w10943w(i) <= wire_cata_12_cordic_atan_w_lg_indexbit10942w(0) AND wire_cata_12_cordic_atan_w_valuenode_12_w_range10941w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_12_cordic_atan_w_lg_indexbit10940w(i) <= indexbit AND wire_cata_12_cordic_atan_w_valuenode_14_w_range10939w(i);
	END GENERATE loop7;
	wire_cata_12_cordic_atan_w_lg_indexbit10942w(0) <= NOT indexbit;
	arctan <= (wire_cata_12_cordic_atan_w_lg_w_lg_indexbit10942w10943w OR wire_cata_12_cordic_atan_w_lg_indexbit10940w);
	valuenode_12_w <= "000000000000001111111111111111111111111010101011";
	valuenode_14_w <= "000000000000000011111111111111111111111111111011";
	wire_cata_12_cordic_atan_w_valuenode_12_w_range10941w <= valuenode_12_w(47 DOWNTO 14);
	wire_cata_12_cordic_atan_w_valuenode_14_w_range10939w <= valuenode_14_w(45 DOWNTO 12);

 END RTL; --sinhw_altfp_sincos_cordic_atan_n6b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=13 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_o6b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_o6b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_o6b IS

	 SIGNAL  wire_cata_13_cordic_atan_w_lg_w_lg_indexbit10948w10949w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_w_lg_indexbit10946w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_w_lg_indexbit10948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_13_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_15_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_w_valuenode_13_w_range10947w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_w_valuenode_15_w_range10945w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop8 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_13_cordic_atan_w_lg_w_lg_indexbit10948w10949w(i) <= wire_cata_13_cordic_atan_w_lg_indexbit10948w(0) AND wire_cata_13_cordic_atan_w_valuenode_13_w_range10947w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_13_cordic_atan_w_lg_indexbit10946w(i) <= indexbit AND wire_cata_13_cordic_atan_w_valuenode_15_w_range10945w(i);
	END GENERATE loop9;
	wire_cata_13_cordic_atan_w_lg_indexbit10948w(0) <= NOT indexbit;
	arctan <= (wire_cata_13_cordic_atan_w_lg_w_lg_indexbit10948w10949w OR wire_cata_13_cordic_atan_w_lg_indexbit10946w);
	valuenode_13_w <= "000000000000000111111111111111111111111111010101";
	valuenode_15_w <= "000000000000000001111111111111111111111111111111";
	wire_cata_13_cordic_atan_w_valuenode_13_w_range10947w <= valuenode_13_w(47 DOWNTO 14);
	wire_cata_13_cordic_atan_w_valuenode_15_w_range10945w <= valuenode_15_w(45 DOWNTO 12);

 END RTL; --sinhw_altfp_sincos_cordic_atan_o6b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=1 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_55b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_55b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_55b IS

	 SIGNAL  wire_cata_1_cordic_atan_w_lg_w_lg_indexbit10954w10955w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_w_lg_indexbit10952w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_w_lg_indexbit10954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_1_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_3_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_w_valuenode_1_w_range10953w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_w_valuenode_3_w_range10951w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop10 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_1_cordic_atan_w_lg_w_lg_indexbit10954w10955w(i) <= wire_cata_1_cordic_atan_w_lg_indexbit10954w(0) AND wire_cata_1_cordic_atan_w_valuenode_1_w_range10953w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_1_cordic_atan_w_lg_indexbit10952w(i) <= indexbit AND wire_cata_1_cordic_atan_w_valuenode_3_w_range10951w(i);
	END GENERATE loop11;
	wire_cata_1_cordic_atan_w_lg_indexbit10954w(0) <= NOT indexbit;
	arctan <= (wire_cata_1_cordic_atan_w_lg_w_lg_indexbit10954w10955w OR wire_cata_1_cordic_atan_w_lg_indexbit10952w);
	valuenode_1_w <= "000111011010110001100111000001010110000110111011";
	valuenode_3_w <= "000001111111010101101110101001101010101100001100";
	wire_cata_1_cordic_atan_w_valuenode_1_w_range10953w <= valuenode_1_w(47 DOWNTO 14);
	wire_cata_1_cordic_atan_w_valuenode_3_w_range10951w <= valuenode_3_w(45 DOWNTO 12);

 END RTL; --sinhw_altfp_sincos_cordic_atan_55b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=2 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_65b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_65b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_65b IS

	 SIGNAL  wire_cata_2_cordic_atan_w_lg_w_lg_indexbit10960w10961w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_w_lg_indexbit10958w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_w_lg_indexbit10960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_2_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_4_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_w_valuenode_2_w_range10959w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_w_valuenode_4_w_range10957w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop12 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_2_cordic_atan_w_lg_w_lg_indexbit10960w10961w(i) <= wire_cata_2_cordic_atan_w_lg_indexbit10960w(0) AND wire_cata_2_cordic_atan_w_valuenode_2_w_range10959w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_2_cordic_atan_w_lg_indexbit10958w(i) <= indexbit AND wire_cata_2_cordic_atan_w_valuenode_4_w_range10957w(i);
	END GENERATE loop13;
	wire_cata_2_cordic_atan_w_lg_indexbit10960w(0) <= NOT indexbit;
	arctan <= (wire_cata_2_cordic_atan_w_lg_w_lg_indexbit10960w10961w OR wire_cata_2_cordic_atan_w_lg_indexbit10958w);
	valuenode_2_w <= "000011111010110110111010111111001001011001000000";
	valuenode_4_w <= "000000111111111010101011011101101110010110100000";
	wire_cata_2_cordic_atan_w_valuenode_2_w_range10959w <= valuenode_2_w(47 DOWNTO 14);
	wire_cata_2_cordic_atan_w_valuenode_4_w_range10957w <= valuenode_4_w(45 DOWNTO 12);

 END RTL; --sinhw_altfp_sincos_cordic_atan_65b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=3 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_75b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_75b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_75b IS

	 SIGNAL  wire_cata_3_cordic_atan_w_lg_w_lg_indexbit10966w10967w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_w_lg_indexbit10964w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_w_lg_indexbit10966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_3_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_5_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_w_valuenode_3_w_range10965w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_w_valuenode_5_w_range10963w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop14 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_3_cordic_atan_w_lg_w_lg_indexbit10966w10967w(i) <= wire_cata_3_cordic_atan_w_lg_indexbit10966w(0) AND wire_cata_3_cordic_atan_w_valuenode_3_w_range10965w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_3_cordic_atan_w_lg_indexbit10964w(i) <= indexbit AND wire_cata_3_cordic_atan_w_valuenode_5_w_range10963w(i);
	END GENERATE loop15;
	wire_cata_3_cordic_atan_w_lg_indexbit10966w(0) <= NOT indexbit;
	arctan <= (wire_cata_3_cordic_atan_w_lg_w_lg_indexbit10966w10967w OR wire_cata_3_cordic_atan_w_lg_indexbit10964w);
	valuenode_3_w <= "000001111111010101101110101001101010101100001100";
	valuenode_5_w <= "000000011111111111010101010110111011101010010111";
	wire_cata_3_cordic_atan_w_valuenode_3_w_range10965w <= valuenode_3_w(47 DOWNTO 14);
	wire_cata_3_cordic_atan_w_valuenode_5_w_range10963w <= valuenode_5_w(45 DOWNTO 12);

 END RTL; --sinhw_altfp_sincos_cordic_atan_75b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=4 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_85b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_85b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_85b IS

	 SIGNAL  wire_cata_4_cordic_atan_w_lg_w_lg_indexbit10972w10973w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_w_lg_indexbit10970w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_w_lg_indexbit10972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_4_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_6_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_w_valuenode_4_w_range10971w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_w_valuenode_6_w_range10969w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop16 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_4_cordic_atan_w_lg_w_lg_indexbit10972w10973w(i) <= wire_cata_4_cordic_atan_w_lg_indexbit10972w(0) AND wire_cata_4_cordic_atan_w_valuenode_4_w_range10971w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_4_cordic_atan_w_lg_indexbit10970w(i) <= indexbit AND wire_cata_4_cordic_atan_w_valuenode_6_w_range10969w(i);
	END GENERATE loop17;
	wire_cata_4_cordic_atan_w_lg_indexbit10972w(0) <= NOT indexbit;
	arctan <= (wire_cata_4_cordic_atan_w_lg_w_lg_indexbit10972w10973w OR wire_cata_4_cordic_atan_w_lg_indexbit10970w);
	valuenode_4_w <= "000000111111111010101011011101101110010110100000";
	valuenode_6_w <= "000000001111111111111010101010101101110111011100";
	wire_cata_4_cordic_atan_w_valuenode_4_w_range10971w <= valuenode_4_w(47 DOWNTO 14);
	wire_cata_4_cordic_atan_w_valuenode_6_w_range10969w <= valuenode_6_w(45 DOWNTO 12);

 END RTL; --sinhw_altfp_sincos_cordic_atan_85b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=5 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_95b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_95b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_95b IS

	 SIGNAL  wire_cata_5_cordic_atan_w_lg_w_lg_indexbit10978w10979w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_w_lg_indexbit10976w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_w_lg_indexbit10978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_5_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_7_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_w_valuenode_5_w_range10977w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_w_valuenode_7_w_range10975w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop18 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_5_cordic_atan_w_lg_w_lg_indexbit10978w10979w(i) <= wire_cata_5_cordic_atan_w_lg_indexbit10978w(0) AND wire_cata_5_cordic_atan_w_valuenode_5_w_range10977w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_5_cordic_atan_w_lg_indexbit10976w(i) <= indexbit AND wire_cata_5_cordic_atan_w_valuenode_7_w_range10975w(i);
	END GENERATE loop19;
	wire_cata_5_cordic_atan_w_lg_indexbit10978w(0) <= NOT indexbit;
	arctan <= (wire_cata_5_cordic_atan_w_lg_w_lg_indexbit10978w10979w OR wire_cata_5_cordic_atan_w_lg_indexbit10976w);
	valuenode_5_w <= "000000011111111111010101010110111011101010010111";
	valuenode_7_w <= "000000000111111111111111010101010101011011101111";
	wire_cata_5_cordic_atan_w_valuenode_5_w_range10977w <= valuenode_5_w(47 DOWNTO 14);
	wire_cata_5_cordic_atan_w_valuenode_7_w_range10975w <= valuenode_7_w(45 DOWNTO 12);

 END RTL; --sinhw_altfp_sincos_cordic_atan_95b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=6 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_a5b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_a5b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_a5b IS

	 SIGNAL  wire_cata_6_cordic_atan_w_lg_w_lg_indexbit10984w10985w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_w_lg_indexbit10982w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_w_lg_indexbit10984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_6_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_8_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_w_valuenode_6_w_range10983w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_w_valuenode_8_w_range10981w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop20 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_6_cordic_atan_w_lg_w_lg_indexbit10984w10985w(i) <= wire_cata_6_cordic_atan_w_lg_indexbit10984w(0) AND wire_cata_6_cordic_atan_w_valuenode_6_w_range10983w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_6_cordic_atan_w_lg_indexbit10982w(i) <= indexbit AND wire_cata_6_cordic_atan_w_valuenode_8_w_range10981w(i);
	END GENERATE loop21;
	wire_cata_6_cordic_atan_w_lg_indexbit10984w(0) <= NOT indexbit;
	arctan <= (wire_cata_6_cordic_atan_w_lg_w_lg_indexbit10984w10985w OR wire_cata_6_cordic_atan_w_lg_indexbit10982w);
	valuenode_6_w <= "000000001111111111111010101010101101110111011100";
	valuenode_8_w <= "000000000011111111111111111010101010101010110111";
	wire_cata_6_cordic_atan_w_valuenode_6_w_range10983w <= valuenode_6_w(47 DOWNTO 14);
	wire_cata_6_cordic_atan_w_valuenode_8_w_range10981w <= valuenode_8_w(45 DOWNTO 12);

 END RTL; --sinhw_altfp_sincos_cordic_atan_a5b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=7 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_b5b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_b5b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_b5b IS

	 SIGNAL  wire_cata_7_cordic_atan_w_lg_w_lg_indexbit10990w10991w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_w_lg_indexbit10988w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_w_lg_indexbit10990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_7_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_9_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_w_valuenode_7_w_range10989w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_w_valuenode_9_w_range10987w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop22 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_7_cordic_atan_w_lg_w_lg_indexbit10990w10991w(i) <= wire_cata_7_cordic_atan_w_lg_indexbit10990w(0) AND wire_cata_7_cordic_atan_w_valuenode_7_w_range10989w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_7_cordic_atan_w_lg_indexbit10988w(i) <= indexbit AND wire_cata_7_cordic_atan_w_valuenode_9_w_range10987w(i);
	END GENERATE loop23;
	wire_cata_7_cordic_atan_w_lg_indexbit10990w(0) <= NOT indexbit;
	arctan <= (wire_cata_7_cordic_atan_w_lg_w_lg_indexbit10990w10991w OR wire_cata_7_cordic_atan_w_lg_indexbit10988w);
	valuenode_7_w <= "000000000111111111111111010101010101011011101111";
	valuenode_9_w <= "000000000001111111111111111111010101010101010110";
	wire_cata_7_cordic_atan_w_valuenode_7_w_range10989w <= valuenode_7_w(47 DOWNTO 14);
	wire_cata_7_cordic_atan_w_valuenode_9_w_range10987w <= valuenode_9_w(45 DOWNTO 12);

 END RTL; --sinhw_altfp_sincos_cordic_atan_b5b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=8 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_c5b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_c5b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_c5b IS

	 SIGNAL  wire_cata_8_cordic_atan_w_lg_w_lg_indexbit10996w10997w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_w_lg_indexbit10994w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_w_lg_indexbit10996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_10_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_8_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_w_valuenode_10_w_range10993w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_w_valuenode_8_w_range10995w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop24 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_8_cordic_atan_w_lg_w_lg_indexbit10996w10997w(i) <= wire_cata_8_cordic_atan_w_lg_indexbit10996w(0) AND wire_cata_8_cordic_atan_w_valuenode_8_w_range10995w(i);
	END GENERATE loop24;
	loop25 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_8_cordic_atan_w_lg_indexbit10994w(i) <= indexbit AND wire_cata_8_cordic_atan_w_valuenode_10_w_range10993w(i);
	END GENERATE loop25;
	wire_cata_8_cordic_atan_w_lg_indexbit10996w(0) <= NOT indexbit;
	arctan <= (wire_cata_8_cordic_atan_w_lg_w_lg_indexbit10996w10997w OR wire_cata_8_cordic_atan_w_lg_indexbit10994w);
	valuenode_10_w <= "000000000000111111111111111111111010101010101011";
	valuenode_8_w <= "000000000011111111111111111010101010101010110111";
	wire_cata_8_cordic_atan_w_valuenode_10_w_range10993w <= valuenode_10_w(45 DOWNTO 12);
	wire_cata_8_cordic_atan_w_valuenode_8_w_range10995w <= valuenode_8_w(47 DOWNTO 14);

 END RTL; --sinhw_altfp_sincos_cordic_atan_c5b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=2 START=9 WIDTH=34 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_atan_d5b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_atan_d5b;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_atan_d5b IS

	 SIGNAL  wire_cata_9_cordic_atan_w_lg_w_lg_indexbit11002w11003w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_w_lg_indexbit11000w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_w_lg_indexbit11002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_11_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_9_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_w_valuenode_11_w_range10999w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_w_valuenode_9_w_range11001w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
 BEGIN

	loop26 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_9_cordic_atan_w_lg_w_lg_indexbit11002w11003w(i) <= wire_cata_9_cordic_atan_w_lg_indexbit11002w(0) AND wire_cata_9_cordic_atan_w_valuenode_9_w_range11001w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 33 GENERATE 
		wire_cata_9_cordic_atan_w_lg_indexbit11000w(i) <= indexbit AND wire_cata_9_cordic_atan_w_valuenode_11_w_range10999w(i);
	END GENERATE loop27;
	wire_cata_9_cordic_atan_w_lg_indexbit11002w(0) <= NOT indexbit;
	arctan <= (wire_cata_9_cordic_atan_w_lg_w_lg_indexbit11002w11003w OR wire_cata_9_cordic_atan_w_lg_indexbit11000w);
	valuenode_11_w <= "000000000000011111111111111111111111010101010101";
	valuenode_9_w <= "000000000001111111111111111111010101010101010110";
	wire_cata_9_cordic_atan_w_valuenode_11_w_range10999w <= valuenode_11_w(45 DOWNTO 12);
	wire_cata_9_cordic_atan_w_valuenode_9_w_range11001w <= valuenode_9_w(47 DOWNTO 14);

 END RTL; --sinhw_altfp_sincos_cordic_atan_d5b


--altfp_sincos_cordic_start CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" WIDTH=34 index value
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_mux 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_start_709 IS 
	 PORT 
	 ( 
		 index	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
		 value	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0)
	 ); 
 END sinhw_altfp_sincos_cordic_start_709;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_start_709 IS

	 SIGNAL  wire_mux1_data	:	STD_LOGIC_VECTOR (543 DOWNTO 0);
	 SIGNAL  wire_mux1_data_2d	:	STD_LOGIC_2D(15 DOWNTO 0, 33 DOWNTO 0);
	 SIGNAL  wire_mux1_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  valuenode_0_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_10_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_11_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_12_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_13_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_14_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_15_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_1_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_2_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_3_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_4_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_5_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_6_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_7_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_8_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_9_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
 BEGIN

	value <= wire_mux1_result;
	valuenode_0_w <= "001001101101110100111011011010100001";
	valuenode_10_w <= "001111111111111111111101010101010101";
	valuenode_11_w <= "001111111111111111111111010101010101";
	valuenode_12_w <= "001111111111111111111111111101010101";
	valuenode_13_w <= "001111111111111111111111110101010101";
	valuenode_14_w <= "001111111111111111111111111111110101";
	valuenode_15_w <= "001111111111111111111111111111010101";
	valuenode_1_w <= "001101101111011001010110110001011010";
	valuenode_2_w <= "001111010111001100011101111111111011";
	valuenode_3_w <= "001111110101011101000011101100100100";
	valuenode_4_w <= "001111111101010101110100100001100000";
	valuenode_5_w <= "001111111111010101010111010010011001";
	valuenode_6_w <= "001111111111110101010101011101001010";
	valuenode_7_w <= "001111111111111101010101010101110101";
	valuenode_8_w <= "001111111111111111010101010101010111";
	valuenode_9_w <= "001111111111111111110101010101010101";
	wire_mux1_data <= ( valuenode_15_w(35 DOWNTO 2) & valuenode_14_w(35 DOWNTO 2) & valuenode_13_w(35 DOWNTO 2) & valuenode_12_w(35 DOWNTO 2) & valuenode_11_w(35 DOWNTO 2) & valuenode_10_w(35 DOWNTO 2) & valuenode_9_w(35 DOWNTO 2) & valuenode_8_w(35 DOWNTO 2) & valuenode_7_w(35 DOWNTO 2) & valuenode_6_w(35 DOWNTO 2) & valuenode_5_w(35 DOWNTO 2) & valuenode_4_w(35 DOWNTO 2) & valuenode_3_w(35 DOWNTO 2) & valuenode_2_w(35 DOWNTO 2) & valuenode_1_w(35 DOWNTO 2) & valuenode_0_w(35 DOWNTO 2));
	loop28 : FOR i IN 0 TO 15 GENERATE
		loop29 : FOR j IN 0 TO 33 GENERATE
			wire_mux1_data_2d(i, j) <= wire_mux1_data(i*34+j);
		END GENERATE loop29;
	END GENERATE loop28;
	mux1 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 16,
		LPM_WIDTH => 34,
		LPM_WIDTHS => 4
	  )
	  PORT MAP ( 
		data => wire_mux1_data_2d,
		result => wire_mux1_result,
		sel => index
	  );

 END RTL; --sinhw_altfp_sincos_cordic_start_709

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 39 lpm_mult 1 lpm_mux 1 reg 1598 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_cordic_m_e5e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 indexbit	:	IN  STD_LOGIC := '0';
		 radians	:	IN  STD_LOGIC_VECTOR (33 DOWNTO 0) := (OTHERS => '0');
		 sincos	:	OUT  STD_LOGIC_VECTOR (33 DOWNTO 0);
		 sincosbit	:	IN  STD_LOGIC := '0'
	 ); 
 END sinhw_altfp_sincos_cordic_m_e5e;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_cordic_m_e5e IS

	 SIGNAL  wire_cata_0_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_arctan	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cxs_value	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL	 cdaff_0	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cdaff_1	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cdaff_2	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 indexbitff	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_indexbitff_w_lg_w_q_range581w679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range610w8590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range613w9392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range616w10189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range10749w10752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range583w1147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range586w1994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range589w2836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range592w3673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range595w4505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range598w5332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range601w6154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range604w6971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range607w7783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range10749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 sincosbitff	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_sincosbitff_w_lg_w_q_range668w10739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sincosbitff_w_lg_w_q_range10746w10747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sincosbitff_w_q_range668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sincosbitff_w_q_range10746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 sincosff	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_0	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range680w681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range721w733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range721w722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range726w738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range726w727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range731w743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range731w732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range736w748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range736w737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range741w753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range741w742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range746w758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range746w747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range751w763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range751w752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range756w768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range756w757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range761w773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range761w762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range766w778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range766w767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range687w688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range771w783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range771w772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range776w788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range776w777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range781w793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range781w782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range786w798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range786w787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range791w803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range791w792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range796w808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range796w797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range801w813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range801w802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range806w818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range806w807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range811w823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range811w812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range816w828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range816w817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range677w693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range677w678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range821w833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range821w822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range826w838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range826w827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range831w841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range831w832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range836w837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range685w698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range685w686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range691w703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range691w692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range696w708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range696w697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range701w713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range701w702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range706w718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range706w707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range711w723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range711w712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range716w728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range716w717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range836w843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range680w681w682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range721w733w734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range726w738w739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range731w743w744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range736w748w749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range741w753w754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range746w758w759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range751w763w764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range756w768w769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range761w773w774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range766w778w779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range687w688w689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range771w783w784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range776w788w789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range781w793w794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range786w798w799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range791w803w804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range796w808w809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range801w813w814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range806w818w819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range811w823w824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range816w828w829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range677w693w694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range821w833w834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range826w838w839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range685w698w699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range691w703w704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range696w708w709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range701w713w714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range706w718w719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range711w723w724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range716w728w729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 x_pipeff_1	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_10	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_11	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_12	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_13	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_x_pipeff_13_w_lg_q10744w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_13_w_lg_q10741w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL	 x_pipeff_2	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_3	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_4	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_5	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_6	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_7	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_8	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_9	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 y_pipeff_0	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 y_pipeff_1	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range913w914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range919w920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range925w926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range931w932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range937w938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range943w944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range949w950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range955w956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range961w962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range967w968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range860w861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range973w974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range979w980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range985w986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range991w992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range997w998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1003w1004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1009w1010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1015w1016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1021w1022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1027w1028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range865w866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1033w1034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1039w1040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range1045w1046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range845w846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range871w872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range877w878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range883w884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range889w890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range895w896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range901w902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range907w908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range1045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_10	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8384w8385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8389w8390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8395w8396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8401w8402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8407w8408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8413w8414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8419w8420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8425w8426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8431w8432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8437w8438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8443w8444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8449w8450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8455w8456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8461w8462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8467w8468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8473w8474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8479w8480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8485w8486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8491w8492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8497w8498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8503w8504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8509w8510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8515w8516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range8333w8334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range8333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_11	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9195w9196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9200w9201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9206w9207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9212w9213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9218w9219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9224w9225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9230w9231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9236w9237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9242w9243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9248w9249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9254w9255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9260w9261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9266w9267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9272w9273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9278w9279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9284w9285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9290w9291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9296w9297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9302w9303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9308w9309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9314w9315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9320w9321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range9140w9141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range9140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_12	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10001w10002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10006w10007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10012w10013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10018w10019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10024w10025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10030w10031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10036w10037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10042w10043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10048w10049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10054w10055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10060w10061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10066w10067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10072w10073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10078w10079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10084w10085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10090w10091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10096w10097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10102w10103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10108w10109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10114w10115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range10120w10121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9942w9943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range10120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_13	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_13_w_lg_q10740w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_13_w_lg_q10743w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL	 y_pipeff_2	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1763w1764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1769w1770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1775w1776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1781w1782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1787w1788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1793w1794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1799w1800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1805w1806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1811w1812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1817w1818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1823w1824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1829w1830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1835w1836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1841w1842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1847w1848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1853w1854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1859w1860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1865w1866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1871w1872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1877w1878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1716w1717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1883w1884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1889w1890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1895w1896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1697w1698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1721w1722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1727w1728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1733w1734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1739w1740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1745w1746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1751w1752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1757w1758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_3	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2608w2609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2614w2615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2620w2621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2626w2627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2632w2633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2638w2639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2644w2645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2650w2651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2656w2657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2662w2663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2668w2669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2674w2675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2680w2681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2686w2687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2692w2693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2698w2699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2704w2705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2710w2711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2716w2717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2722w2723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2728w2729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2734w2735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2740w2741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2544w2545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2567w2568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2572w2573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2578w2579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2584w2585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2590w2591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2596w2597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2602w2603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_4	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3448w3449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3454w3455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3460w3461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3466w3467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3472w3473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3478w3479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3484w3485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3490w3491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3496w3497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3502w3503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3508w3509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3514w3515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3520w3521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3526w3527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3532w3533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3538w3539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3544w3545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3550w3551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3556w3557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3562w3563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3568w3569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3574w3575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3580w3581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3386w3387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3413w3414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3418w3419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3424w3425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3430w3431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3436w3437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3442w3443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_5	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4283w4284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4289w4290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4295w4296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4301w4302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4307w4308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4313w4314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4319w4320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4325w4326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4331w4332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4337w4338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4343w4344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4349w4350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4355w4356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4361w4362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4367w4368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4373w4374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4379w4380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4385w4386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4391w4392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4397w4398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4403w4404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4409w4410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4415w4416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4223w4224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4254w4255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4259w4260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4265w4266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4271w4272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4277w4278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_6	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5113w5114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5119w5120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5125w5126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5131w5132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5137w5138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5143w5144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5149w5150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5155w5156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5161w5162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5167w5168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5173w5174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5179w5180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5185w5186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5191w5192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5197w5198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5203w5204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5209w5210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5215w5216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5221w5222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5227w5228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5233w5234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5239w5240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5245w5246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5055w5056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5090w5091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5095w5096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5101w5102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range5107w5108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range5107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_7	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5938w5939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5944w5945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5950w5951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5956w5957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5962w5963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5968w5969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5974w5975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5980w5981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5986w5987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5992w5993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5998w5999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6004w6005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6010w6011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6016w6017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6022w6023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6028w6029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6034w6035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6040w6041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6046w6047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6052w6053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6058w6059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6064w6065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range6070w6071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5882w5883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5921w5922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5926w5927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5932w5933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range6070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_8	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6758w6759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6764w6765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6770w6771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6776w6777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6782w6783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6788w6789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6794w6795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6800w6801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6806w6807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6812w6813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6818w6819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6824w6825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6830w6831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6836w6837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6842w6843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6848w6849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6854w6855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6860w6861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6866w6867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6872w6873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6878w6879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6884w6885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6890w6891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6704w6705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6747w6748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6752w6753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_9	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7573w7574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7579w7580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7585w7586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7591w7592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7597w7598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7603w7604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7609w7610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7615w7616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7621w7622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7627w7628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7633w7634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7639w7640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7645w7646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7651w7652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7657w7658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7663w7664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7669w7670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7675w7676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7681w7682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7687w7688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7693w7694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7699w7700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7705w7706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7521w7522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7568w7569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_0	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 z_pipeff_1	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_1_w_q_range1421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_10	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_10_w_q_range8864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_11	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_11_w_q_range9666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_12	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_12_w_q_range10463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_13	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 z_pipeff_2	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_2_w_q_range2268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_3	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_3_w_q_range3110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_4	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_4_w_q_range3947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_5	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_5_w_q_range4779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_6	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_6_w_q_range5606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_7	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_7_w_q_range6428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_8	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_8_w_q_range7245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_9	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_9_w_q_range8057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sincos_add_cin	:	STD_LOGIC;
	 SIGNAL  wire_sincos_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_10_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_11_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_12_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_13_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_2_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_3_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_4_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_5_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_6_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_7_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_8_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_9_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipeff1_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_10_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_11_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_12_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_13_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_2_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_3_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_4_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_5_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_6_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_7_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_8_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_9_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipeff1_sub_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_10_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_11_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_12_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_13_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_2_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_3_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_4_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_5_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_6_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_7_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_8_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_9_add_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_cmx_result	:	STD_LOGIC_VECTOR (67 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_indexpointnum_w409w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10753w10754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10794w10806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10794w10795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10799w10811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10799w10800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10804w10816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10804w10805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10809w10821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10809w10810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10814w10826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10814w10815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10819w10831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10819w10820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10824w10836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10824w10825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10829w10841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10829w10830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10834w10846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10834w10835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10839w10851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10839w10840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10760w10761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10844w10856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10844w10845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10849w10861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10849w10850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10854w10866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10854w10855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10859w10871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10859w10860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10864w10876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10864w10865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10869w10881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10869w10870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10874w10886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10874w10875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10879w10891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10879w10880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10884w10896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10884w10885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10889w10901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10889w10890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10750w10766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10750w10751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10894w10906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10894w10895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10899w10911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10899w10900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10904w10914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10904w10905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10758w10771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10758w10759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10764w10776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10764w10765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10769w10781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10769w10770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10774w10786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10774w10775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10779w10791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10779w10780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10784w10796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10784w10785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10789w10801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10789w10790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range410w413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range410w420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range458w461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range458w470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range463w466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range463w475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range468w471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range468w480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range473w476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range473w485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range478w481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range478w490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range483w486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range483w495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range488w491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range488w500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range493w496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range493w505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range498w501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range498w510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range503w506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range503w515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range415w417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range415w425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range508w511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range508w520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range513w516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range513w525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range518w521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range518w530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range523w526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range523w535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range528w531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range528w540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range533w536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range533w545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range538w541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range538w550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range543w546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range543w555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range548w551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range548w560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range553w556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range553w565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range418w421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range418w430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range558w561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range558w570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range563w566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range563w575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range568w571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range573w576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range423w426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range423w435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range428w431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range428w440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range433w436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range433w445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range438w441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range438w450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range443w446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range443w455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range448w451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range448w460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range453w456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range453w465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7570w7784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7629w7866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7635w7874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7641w7882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7647w7890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7653w7898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7659w7906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7665w7914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7671w7922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7677w7930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7683w7938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7575w7794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7689w7946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7695w7954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7701w7962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7707w7970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7711w7978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7523w7986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7528w7994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7530w8002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7532w8010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7534w8018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7581w7802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7536w8026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7538w8034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7540w8042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7542w8050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7587w7810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7593w7818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7599w7826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7605w7834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7611w7842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7617w7850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7623w7858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8386w8591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8445w8673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8451w8681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8457w8689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8463w8697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8469w8705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8475w8713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8481w8721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8487w8729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8493w8737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8499w8745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8391w8601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8505w8753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8511w8761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8517w8769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8521w8777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8335w8785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8340w8793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8342w8801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8344w8809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8346w8817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8348w8825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8397w8609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8350w8833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8352w8841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8354w8849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8356w8857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8403w8617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8409w8625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8415w8633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8421w8641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8427w8649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8433w8657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8439w8665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9197w9393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9256w9475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9262w9483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9268w9491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9274w9499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9280w9507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9286w9515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9292w9523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9298w9531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9304w9539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9310w9547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9202w9403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9316w9555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9322w9563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9326w9571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9142w9579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9147w9587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9149w9595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9151w9603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9153w9611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9155w9619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9157w9627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9208w9411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9159w9635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9161w9643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9163w9651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9165w9659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9214w9419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9220w9427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9226w9435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9232w9443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9238w9451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9244w9459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9250w9467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10003w10190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10062w10272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10068w10280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10074w10288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10080w10296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10086w10304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10092w10312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10098w10320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10104w10328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10110w10336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10116w10344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10008w10200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10122w10352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10126w10360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9944w10368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9949w10376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9951w10384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9953w10392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9955w10400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9957w10408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9959w10416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9961w10424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10014w10208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9963w10432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9965w10440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9967w10448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9969w10456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10020w10216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10026w10224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10032w10232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10038w10240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10044w10248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10050w10256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10056w10264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range862w1148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range921w1230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range927w1238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range933w1246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range939w1254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range945w1262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range951w1270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range957w1278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range963w1286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range969w1294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range975w1302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range867w1158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range981w1310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range987w1318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range993w1326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range999w1334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1005w1342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1011w1350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1017w1358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1023w1366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1029w1374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1035w1382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range873w1166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1041w1390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1047w1398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1051w1406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range847w1414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range879w1174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range885w1182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range891w1190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range897w1198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range903w1206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range909w1214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range915w1222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1718w1995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1777w2077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1783w2085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1789w2093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1795w2101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1801w2109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1807w2117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1813w2125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1819w2133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1825w2141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1831w2149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1723w2005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1837w2157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1843w2165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1849w2173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1855w2181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1861w2189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1867w2197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1873w2205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1879w2213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1885w2221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1891w2229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1729w2013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1897w2237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1901w2245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1699w2253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1704w2261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1735w2021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1741w2029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1747w2037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1753w2045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1759w2053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1765w2061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1771w2069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2569w2837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2628w2919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2634w2927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2640w2935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2646w2943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2652w2951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2658w2959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2664w2967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2670w2975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2676w2983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2682w2991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2574w2847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2688w2999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2694w3007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2700w3015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2706w3023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2712w3031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2718w3039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2724w3047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2730w3055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2736w3063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2742w3071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2580w2855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2746w3079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2546w3087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2551w3095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2553w3103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2586w2863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2592w2871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2598w2879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2604w2887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2610w2895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2616w2903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2622w2911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3415w3674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3474w3756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3480w3764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3486w3772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3492w3780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3498w3788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3504w3796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3510w3804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3516w3812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3522w3820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3528w3828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3420w3684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3534w3836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3540w3844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3546w3852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3552w3860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3558w3868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3564w3876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3570w3884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3576w3892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3582w3900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3586w3908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3426w3692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3388w3916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3393w3924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3395w3932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3397w3940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3432w3700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3438w3708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3444w3716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3450w3724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3456w3732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3462w3740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3468w3748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4256w4506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4315w4588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4321w4596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4327w4604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4333w4612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4339w4620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4345w4628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4351w4636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4357w4644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4363w4652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4369w4660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4261w4516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4375w4668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4381w4676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4387w4684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4393w4692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4399w4700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4405w4708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4411w4716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4417w4724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4421w4732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4225w4740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4267w4524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4230w4748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4232w4756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4234w4764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4236w4772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4273w4532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4279w4540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4285w4548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4291w4556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4297w4564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4303w4572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4309w4580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5092w5333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5151w5415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5157w5423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5163w5431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5169w5439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5175w5447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5181w5455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5187w5463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5193w5471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5199w5479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5205w5487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5097w5343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5211w5495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5217w5503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5223w5511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5229w5519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5235w5527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5241w5535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5247w5543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5251w5551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5057w5559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5062w5567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5103w5351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5064w5575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5066w5583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5068w5591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5070w5599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5109w5359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5115w5367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5121w5375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5127w5383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5133w5391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5139w5399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5145w5407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5923w6155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5982w6237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5988w6245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5994w6253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6000w6261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6006w6269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6012w6277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6018w6285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6024w6293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6030w6301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6036w6309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5928w6165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6042w6317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6048w6325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6054w6333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6060w6341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6066w6349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6072w6357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6076w6365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5884w6373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5889w6381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5891w6389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5934w6173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5893w6397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5895w6405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5897w6413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5899w6421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5940w6181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5946w6189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5952w6197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5958w6205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5964w6213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5970w6221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5976w6229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6749w6972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6808w7054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6814w7062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6820w7070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6826w7078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6832w7086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6838w7094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6844w7102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6850w7110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6856w7118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6862w7126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6754w6982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6868w7134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6874w7142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6880w7150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6886w7158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6892w7166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6896w7174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6706w7182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6711w7190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6713w7198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6715w7206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6760w6990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6717w7214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6719w7222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6721w7230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6723w7238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6766w6998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6772w7006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6778w7014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6784w7022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6790w7030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6796w7038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6802w7046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7714w7782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7743w7865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7746w7873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7749w7881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7752w7889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7755w7897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7758w7905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7761w7913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7764w7921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7767w7929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7770w7937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7716w7793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7773w7945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7776w7953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7779w7961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7544w7969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7548w7977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7550w7985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7552w7993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7554w8001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7556w8009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7558w8017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7719w7801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7560w8025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7562w8033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7564w8041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7566w8049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7722w7809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7725w7817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7728w7825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7731w7833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7734w7841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7737w7849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7740w7857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8524w8589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8553w8672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8556w8680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8559w8688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8562w8696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8565w8704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8568w8712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8571w8720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8574w8728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8577w8736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8580w8744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8526w8600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8583w8752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8586w8760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8358w8768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8362w8776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8364w8784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8366w8792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8368w8800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8370w8808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8372w8816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8374w8824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8529w8608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8376w8832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8378w8840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8380w8848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8382w8856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8532w8616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8535w8624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8538w8632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8541w8640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8544w8648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8547w8656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8550w8664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9329w9391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9358w9474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9361w9482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9364w9490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9367w9498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9370w9506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9373w9514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9376w9522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9379w9530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9382w9538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9385w9546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9331w9402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9388w9554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9167w9562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9171w9570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9173w9578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9175w9586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9177w9594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9179w9602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9181w9610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9183w9618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9185w9626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9334w9410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9187w9634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9189w9642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9191w9650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9193w9658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9337w9418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9340w9426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9343w9434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9346w9442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9349w9450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9352w9458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9355w9466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10129w10188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10158w10271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10161w10279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10164w10287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10167w10295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10170w10303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10173w10311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10176w10319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10179w10327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10182w10335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10185w10343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10131w10199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9971w10351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9975w10359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9977w10367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9979w10375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9981w10383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9983w10391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9985w10399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9987w10407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9989w10415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9991w10423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10134w10207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9993w10431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9995w10439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9997w10447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9999w10455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10137w10215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10140w10223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10143w10231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10146w10239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10149w10247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10152w10255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10155w10263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1054w1146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1083w1229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1086w1237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1089w1245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1092w1253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1095w1261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1098w1269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1101w1277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1104w1285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1107w1293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1110w1301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1056w1157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1113w1309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1116w1317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1119w1325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1122w1333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1125w1341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1128w1349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1131w1357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1134w1365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1137w1373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1140w1381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1059w1165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1143w1389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range852w1397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range856w1405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range858w1413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1062w1173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1065w1181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1068w1189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1071w1197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1074w1205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1077w1213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1080w1221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1904w1993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1933w2076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1936w2084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1939w2092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1942w2100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1945w2108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1948w2116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1951w2124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1954w2132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1957w2140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1960w2148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1906w2004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1963w2156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1966w2164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1969w2172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1972w2180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1975w2188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1978w2196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1981w2204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1984w2212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1987w2220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1990w2228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1909w2012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1706w2236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1710w2244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1712w2252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1714w2260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1912w2020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1915w2028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1918w2036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1921w2044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1924w2052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1927w2060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1930w2068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2749w2835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2778w2918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2781w2926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2784w2934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2787w2942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2790w2950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2793w2958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2796w2966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2799w2974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2802w2982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2805w2990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2751w2846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2808w2998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2811w3006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2814w3014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2817w3022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2820w3030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2823w3038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2826w3046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2829w3054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2832w3062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2555w3070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2754w2854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2559w3078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2561w3086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2563w3094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2565w3102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2757w2862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2760w2870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2763w2878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2766w2886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2769w2894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2772w2902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2775w2910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3589w3672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3618w3755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3621w3763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3624w3771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3627w3779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3630w3787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3633w3795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3636w3803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3639w3811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3642w3819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3645w3827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3591w3683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3648w3835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3651w3843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3654w3851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3657w3859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3660w3867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3663w3875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3666w3883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3669w3891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3399w3899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3403w3907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3594w3691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3405w3915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3407w3923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3409w3931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3411w3939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3597w3699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3600w3707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3603w3715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3606w3723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3609w3731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3612w3739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3615w3747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4424w4504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4453w4587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4456w4595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4459w4603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4462w4611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4465w4619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4468w4627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4471w4635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4474w4643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4477w4651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4480w4659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4426w4515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4483w4667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4486w4675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4489w4683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4492w4691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4495w4699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4498w4707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4501w4715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4238w4723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4242w4731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4244w4739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4429w4523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4246w4747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4248w4755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4250w4763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4252w4771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4432w4531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4435w4539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4438w4547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4441w4555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4444w4563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4447w4571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4450w4579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5254w5331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5283w5414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5286w5422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5289w5430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5292w5438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5295w5446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5298w5454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5301w5462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5304w5470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5307w5478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5310w5486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5256w5342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5313w5494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5316w5502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5319w5510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5322w5518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5325w5526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5328w5534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5072w5542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5076w5550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5078w5558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5080w5566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5259w5350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5082w5574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5084w5582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5086w5590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5088w5598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5262w5358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5265w5366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5268w5374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5271w5382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5274w5390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5277w5398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5280w5406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6079w6153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6108w6236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6111w6244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6114w6252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6117w6260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6120w6268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6123w6276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6126w6284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6129w6292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6132w6300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6135w6308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6081w6164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6138w6316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6141w6324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6144w6332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6147w6340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6150w6348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5901w6356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5905w6364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5907w6372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5909w6380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5911w6388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6084w6172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5913w6396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5915w6404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5917w6412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5919w6420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6087w6180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6090w6188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6093w6196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6096w6204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6099w6212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6102w6220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6105w6228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6899w6970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6928w7053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6931w7061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6934w7069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6937w7077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6940w7085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6943w7093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6946w7101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6949w7109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6952w7117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6955w7125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6901w6981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6958w7133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6961w7141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6964w7149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6967w7157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6725w7165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6729w7173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6731w7181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6733w7189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6735w7197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6737w7205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6904w6989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6739w7213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6741w7221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6743w7229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6745w7237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6907w6997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6910w7005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6913w7013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6916w7021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6919w7029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6922w7037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6925w7045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7572w7789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7631w7870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7637w7878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7643w7886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7649w7894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7655w7902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7661w7910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7667w7918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7673w7926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7679w7934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7685w7942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7577w7798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7691w7950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7697w7958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7703w7966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7709w7974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7712w7982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7526w7990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7529w7998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7531w8006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7533w8014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7535w8022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7583w7806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7537w8030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7539w8038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7541w8046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7543w8054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7589w7814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7595w7822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7601w7830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7607w7838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7613w7846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7619w7854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7625w7862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8388w8596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8447w8677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8453w8685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8459w8693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8465w8701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8471w8709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8477w8717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8483w8725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8489w8733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8495w8741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8501w8749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8393w8605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8507w8757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8513w8765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8519w8773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8522w8781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8338w8789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8341w8797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8343w8805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8345w8813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8347w8821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8349w8829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8399w8613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8351w8837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8353w8845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8355w8853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8357w8861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8405w8621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8411w8629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8417w8637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8423w8645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8429w8653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8435w8661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8441w8669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9199w9398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9258w9479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9264w9487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9270w9495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9276w9503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9282w9511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9288w9519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9294w9527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9300w9535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9306w9543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9312w9551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9204w9407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9318w9559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9324w9567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9327w9575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9145w9583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9148w9591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9150w9599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9152w9607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9154w9615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9156w9623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9158w9631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9210w9415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9160w9639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9162w9647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9164w9655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9166w9663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9216w9423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9222w9431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9228w9439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9234w9447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9240w9455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9246w9463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9252w9471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10005w10195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10064w10276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10070w10284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10076w10292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10082w10300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10088w10308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10094w10316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10100w10324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10106w10332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10112w10340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10118w10348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10010w10204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10124w10356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10127w10364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9947w10372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9950w10380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9952w10388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9954w10396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9956w10404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9958w10412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9960w10420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9962w10428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10016w10212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9964w10436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9966w10444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9968w10452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9970w10460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10022w10220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10028w10228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10034w10236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10040w10244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10046w10252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10052w10260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10058w10268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range864w1153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range923w1234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range929w1242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range935w1250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range941w1258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range947w1266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range953w1274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range959w1282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range965w1290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range971w1298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range977w1306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range869w1162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range983w1314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range989w1322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range995w1330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1001w1338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1007w1346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1013w1354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1019w1362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1025w1370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1031w1378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1037w1386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range875w1170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1043w1394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1049w1402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1052w1410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range850w1418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range881w1178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range887w1186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range893w1194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range899w1202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range905w1210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range911w1218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range917w1226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1720w2000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1779w2081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1785w2089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1791w2097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1797w2105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1803w2113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1809w2121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1815w2129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1821w2137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1827w2145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1833w2153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1725w2009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1839w2161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1845w2169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1851w2177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1857w2185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1863w2193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1869w2201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1875w2209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1881w2217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1887w2225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1893w2233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1731w2017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1899w2241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1902w2249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1702w2257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1705w2265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1737w2025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1743w2033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1749w2041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1755w2049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1761w2057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1767w2065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1773w2073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2571w2842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2630w2923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2636w2931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2642w2939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2648w2947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2654w2955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2660w2963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2666w2971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2672w2979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2678w2987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2684w2995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2576w2851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2690w3003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2696w3011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2702w3019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2708w3027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2714w3035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2720w3043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2726w3051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2732w3059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2738w3067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2744w3075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2582w2859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2747w3083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2549w3091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2552w3099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2554w3107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2588w2867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2594w2875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2600w2883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2606w2891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2612w2899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2618w2907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2624w2915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3417w3679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3476w3760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3482w3768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3488w3776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3494w3784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3500w3792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3506w3800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3512w3808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3518w3816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3524w3824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3530w3832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3422w3688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3536w3840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3542w3848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3548w3856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3554w3864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3560w3872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3566w3880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3572w3888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3578w3896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3584w3904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3587w3912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3428w3696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3391w3920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3394w3928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3396w3936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3398w3944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3434w3704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3440w3712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3446w3720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3452w3728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3458w3736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3464w3744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3470w3752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4258w4511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4317w4592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4323w4600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4329w4608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4335w4616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4341w4624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4347w4632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4353w4640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4359w4648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4365w4656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4371w4664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4263w4520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4377w4672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4383w4680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4389w4688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4395w4696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4401w4704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4407w4712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4413w4720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4419w4728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4422w4736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4228w4744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4269w4528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4231w4752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4233w4760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4235w4768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4237w4776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4275w4536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4281w4544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4287w4552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4293w4560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4299w4568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4305w4576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4311w4584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5094w5338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5153w5419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5159w5427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5165w5435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5171w5443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5177w5451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5183w5459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5189w5467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5195w5475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5201w5483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5207w5491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5099w5347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5213w5499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5219w5507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5225w5515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5231w5523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5237w5531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5243w5539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5249w5547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5252w5555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5060w5563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5063w5571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5105w5355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5065w5579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5067w5587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5069w5595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5071w5603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5111w5363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5117w5371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5123w5379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5129w5387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5135w5395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5141w5403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5147w5411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5925w6160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5984w6241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5990w6249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5996w6257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6002w6265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6008w6273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6014w6281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6020w6289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6026w6297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6032w6305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6038w6313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5930w6169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6044w6321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6050w6329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6056w6337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6062w6345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6068w6353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6074w6361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6077w6369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5887w6377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5890w6385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5892w6393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5936w6177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5894w6401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5896w6409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5898w6417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5900w6425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5942w6185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5948w6193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5954w6201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5960w6209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5966w6217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5972w6225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5978w6233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6751w6977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6810w7058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6816w7066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6822w7074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6828w7082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6834w7090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6840w7098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6846w7106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6852w7114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6858w7122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6864w7130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6756w6986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6870w7138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6876w7146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6882w7154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6888w7162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6894w7170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6897w7178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6709w7186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6712w7194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6714w7202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6716w7210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6762w6994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6718w7218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6720w7226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6722w7234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6724w7242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6768w7002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6774w7010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6780w7018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6786w7026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6792w7034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6798w7042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6804w7050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7715w7788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7744w7869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7747w7877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7750w7885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7753w7893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7756w7901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7759w7909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7762w7917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7765w7925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7768w7933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7771w7941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7717w7797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7774w7949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7777w7957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7780w7965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7546w7973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7549w7981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7551w7989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7553w7997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7555w8005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7557w8013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7559w8021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7720w7805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7561w8029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7563w8037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7565w8045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7567w8053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7723w7813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7726w7821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7729w7829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7732w7837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7735w7845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7738w7853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7741w7861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8525w8595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8554w8676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8557w8684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8560w8692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8563w8700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8566w8708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8569w8716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8572w8724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8575w8732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8578w8740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8581w8748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8527w8604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8584w8756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8587w8764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8360w8772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8363w8780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8365w8788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8367w8796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8369w8804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8371w8812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8373w8820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8375w8828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8530w8612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8377w8836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8379w8844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8381w8852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8383w8860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8533w8620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8536w8628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8539w8636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8542w8644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8545w8652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8548w8660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8551w8668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9330w9397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9359w9478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9362w9486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9365w9494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9368w9502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9371w9510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9374w9518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9377w9526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9380w9534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9383w9542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9386w9550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9332w9406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9389w9558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9169w9566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9172w9574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9174w9582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9176w9590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9178w9598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9180w9606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9182w9614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9184w9622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9186w9630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9335w9414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9188w9638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9190w9646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9192w9654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9194w9662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9338w9422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9341w9430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9344w9438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9347w9446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9350w9454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9353w9462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9356w9470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10130w10194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10159w10275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10162w10283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10165w10291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10168w10299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10171w10307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10174w10315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10177w10323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10180w10331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10183w10339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10186w10347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10132w10203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9973w10355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9976w10363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9978w10371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9980w10379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9982w10387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9984w10395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9986w10403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9988w10411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9990w10419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9992w10427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10135w10211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9994w10435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9996w10443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9998w10451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10000w10459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10138w10219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10141w10227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10144w10235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10147w10243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10150w10251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10153w10259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10156w10267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1055w1152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1084w1233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1087w1241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1090w1249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1093w1257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1096w1265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1099w1273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1102w1281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1105w1289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1108w1297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1111w1305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1057w1161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1114w1313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1117w1321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1120w1329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1123w1337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1126w1345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1129w1353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1132w1361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1135w1369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1138w1377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1141w1385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1060w1169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1144w1393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range854w1401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range857w1409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range859w1417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1063w1177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1066w1185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1069w1193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1072w1201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1075w1209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1078w1217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1081w1225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1905w1999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1934w2080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1937w2088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1940w2096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1943w2104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1946w2112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1949w2120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1952w2128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1955w2136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1958w2144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1961w2152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1907w2008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1964w2160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1967w2168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1970w2176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1973w2184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1976w2192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1979w2200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1982w2208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1985w2216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1988w2224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1991w2232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1910w2016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1708w2240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1711w2248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1713w2256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1715w2264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1913w2024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1916w2032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1919w2040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1922w2048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1925w2056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1928w2064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1931w2072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2750w2841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2779w2922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2782w2930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2785w2938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2788w2946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2791w2954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2794w2962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2797w2970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2800w2978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2803w2986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2806w2994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2752w2850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2809w3002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2812w3010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2815w3018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2818w3026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2821w3034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2824w3042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2827w3050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2830w3058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2833w3066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2557w3074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2755w2858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2560w3082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2562w3090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2564w3098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2566w3106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2758w2866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2761w2874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2764w2882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2767w2890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2770w2898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2773w2906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2776w2914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3590w3678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3619w3759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3622w3767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3625w3775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3628w3783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3631w3791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3634w3799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3637w3807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3640w3815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3643w3823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3646w3831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3592w3687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3649w3839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3652w3847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3655w3855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3658w3863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3661w3871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3664w3879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3667w3887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3670w3895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3401w3903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3404w3911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3595w3695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3406w3919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3408w3927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3410w3935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3412w3943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3598w3703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3601w3711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3604w3719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3607w3727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3610w3735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3613w3743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3616w3751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4425w4510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4454w4591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4457w4599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4460w4607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4463w4615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4466w4623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4469w4631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4472w4639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4475w4647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4478w4655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4481w4663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4427w4519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4484w4671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4487w4679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4490w4687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4493w4695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4496w4703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4499w4711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4502w4719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4240w4727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4243w4735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4245w4743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4430w4527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4247w4751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4249w4759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4251w4767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4253w4775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4433w4535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4436w4543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4439w4551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4442w4559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4445w4567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4448w4575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4451w4583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5255w5337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5284w5418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5287w5426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5290w5434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5293w5442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5296w5450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5299w5458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5302w5466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5305w5474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5308w5482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5311w5490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5257w5346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5314w5498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5317w5506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5320w5514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5323w5522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5326w5530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5329w5538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5074w5546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5077w5554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5079w5562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5081w5570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5260w5354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5083w5578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5085w5586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5087w5594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5089w5602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5263w5362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5266w5370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5269w5378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5272w5386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5275w5394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5278w5402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5281w5410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6080w6159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6109w6240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6112w6248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6115w6256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6118w6264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6121w6272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6124w6280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6127w6288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6130w6296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6133w6304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6136w6312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6082w6168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6139w6320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6142w6328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6145w6336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6148w6344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6151w6352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5903w6360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5906w6368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5908w6376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5910w6384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5912w6392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6085w6176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5914w6400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5916w6408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5918w6416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5920w6424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6088w6184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6091w6192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6094w6200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6097w6208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6100w6216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6103w6224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6106w6232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6900w6976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6929w7057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6932w7065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6935w7073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6938w7081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6941w7089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6944w7097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6947w7105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6950w7113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6953w7121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6956w7129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6902w6985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6959w7137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6962w7145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6965w7153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6968w7161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6727w7169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6730w7177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6732w7185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6734w7193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6736w7201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6738w7209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6905w6993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6740w7217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6742w7225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6744w7233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6746w7241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6908w7001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6911w7009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6914w7017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6917w7025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6920w7033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6923w7041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6926w7049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_indexbit412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8871w8872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8952w8953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8960w8961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8968w8969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8976w8977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8984w8985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8992w8993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9000w9001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9008w9009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9016w9017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9024w9025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8880w8881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9032w9033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9040w9041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9048w9049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9056w9057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9064w9065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9072w9073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9080w9081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9088w9089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9096w9097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9104w9105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8888w8889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9112w9113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9120w9121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9128w9129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9136w9137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8896w8897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8904w8905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8912w8913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8920w8921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8928w8929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8936w8937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8944w8945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9673w9674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9754w9755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9762w9763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9770w9771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9778w9779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9786w9787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9794w9795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9802w9803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9810w9811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9818w9819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9826w9827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9682w9683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9834w9835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9842w9843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9850w9851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9858w9859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9866w9867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9874w9875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9882w9883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9890w9891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9898w9899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9906w9907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9690w9691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9914w9915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9922w9923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9930w9931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9938w9939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9698w9699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9706w9707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9714w9715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9722w9723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9730w9731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9738w9739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9746w9747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10470w10471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10551w10552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10559w10560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10567w10568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10575w10576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10583w10584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10591w10592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10599w10600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10607w10608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10615w10616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10623w10624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10479w10480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10631w10632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10639w10640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10647w10648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10655w10656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10663w10664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10671w10672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10679w10680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10687w10688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10695w10696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10703w10704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10487w10488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10711w10712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10719w10720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10727w10728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10735w10736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10495w10496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10503w10504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10511w10512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10519w10520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10527w10528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10535w10536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10543w10544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1428w1429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1509w1510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1517w1518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1525w1526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1533w1534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1541w1542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1549w1550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1557w1558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1565w1566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1573w1574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1581w1582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1437w1438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1589w1590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1597w1598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1605w1606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1613w1614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1621w1622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1629w1630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1637w1638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1645w1646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1653w1654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1661w1662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1445w1446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1669w1670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1677w1678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1685w1686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1693w1694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1453w1454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1461w1462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1469w1470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1477w1478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1485w1486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1493w1494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1501w1502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2275w2276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2356w2357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2364w2365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2372w2373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2380w2381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2388w2389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2396w2397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2404w2405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2412w2413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2420w2421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2428w2429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2284w2285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2436w2437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2444w2445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2452w2453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2460w2461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2468w2469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2476w2477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2484w2485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2492w2493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2500w2501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2508w2509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2292w2293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2516w2517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2524w2525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2532w2533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2540w2541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2300w2301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2308w2309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2316w2317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2324w2325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2332w2333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2340w2341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2348w2349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3117w3118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3198w3199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3206w3207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3214w3215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3222w3223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3230w3231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3238w3239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3246w3247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3254w3255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3262w3263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3270w3271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3126w3127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3278w3279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3286w3287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3294w3295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3302w3303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3310w3311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3318w3319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3326w3327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3334w3335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3342w3343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3350w3351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3134w3135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3358w3359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3366w3367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3374w3375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3382w3383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3142w3143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3150w3151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3158w3159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3166w3167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3174w3175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3182w3183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3190w3191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3954w3955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4035w4036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4043w4044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4051w4052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4059w4060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4067w4068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4075w4076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4083w4084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4091w4092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4099w4100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4107w4108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3963w3964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4115w4116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4123w4124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4131w4132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4139w4140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4147w4148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4155w4156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4163w4164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4171w4172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4179w4180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4187w4188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3971w3972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4195w4196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4203w4204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4211w4212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4219w4220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3979w3980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3987w3988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3995w3996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4003w4004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4011w4012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4019w4020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4027w4028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4786w4787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4867w4868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4875w4876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4883w4884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4891w4892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4899w4900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4907w4908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4915w4916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4923w4924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4931w4932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4939w4940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4795w4796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4947w4948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4955w4956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4963w4964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4971w4972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4979w4980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4987w4988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4995w4996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5003w5004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5011w5012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5019w5020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4803w4804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5027w5028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5035w5036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5043w5044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5051w5052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4811w4812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4819w4820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4827w4828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4835w4836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4843w4844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4851w4852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4859w4860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5613w5614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5694w5695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5702w5703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5710w5711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5718w5719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5726w5727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5734w5735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5742w5743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5750w5751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5758w5759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5766w5767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5622w5623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5774w5775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5782w5783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5790w5791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5798w5799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5806w5807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5814w5815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5822w5823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5830w5831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5838w5839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5846w5847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5630w5631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5854w5855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5862w5863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5870w5871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5878w5879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5638w5639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5646w5647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5654w5655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5662w5663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5670w5671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5678w5679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5686w5687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6435w6436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6516w6517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6524w6525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6532w6533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6540w6541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6548w6549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6556w6557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6564w6565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6572w6573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6580w6581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6588w6589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6444w6445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6596w6597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6604w6605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6612w6613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6620w6621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6628w6629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6636w6637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6644w6645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6652w6653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6660w6661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6668w6669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6452w6453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6676w6677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6684w6685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6692w6693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6700w6701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6460w6461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6468w6469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6476w6477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6484w6485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6492w6493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6500w6501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6508w6509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7252w7253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7333w7334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7341w7342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7349w7350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7357w7358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7365w7366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7373w7374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7381w7382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7389w7390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7397w7398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7405w7406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7261w7262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7413w7414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7421w7422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7429w7430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7437w7438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7445w7446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7453w7454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7461w7462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7469w7470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7477w7478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7485w7486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7269w7270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7493w7494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7501w7502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7509w7510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7517w7518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7277w7278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7285w7286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7293w7294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7301w7302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7309w7310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7317w7318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7325w7326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8064w8065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8145w8146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8153w8154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8161w8162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8169w8170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8177w8178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8185w8186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8193w8194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8201w8202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8209w8210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8217w8218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8073w8074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8225w8226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8233w8234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8241w8242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8249w8250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8257w8258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8265w8266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8273w8274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8281w8282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8289w8290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8297w8298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8081w8082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8305w8306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8313w8314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8321w8322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8329w8330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8089w8090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8097w8098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8105w8106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8113w8114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8121w8122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8129w8130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8137w8138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10753w10754w10755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10794w10806w10807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10799w10811w10812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10804w10816w10817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10809w10821w10822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10814w10826w10827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10819w10831w10832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10824w10836w10837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10829w10841w10842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10834w10846w10847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10839w10851w10852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10760w10761w10762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10844w10856w10857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10849w10861w10862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10854w10866w10867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10859w10871w10872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10864w10876w10877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10869w10881w10882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10874w10886w10887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10879w10891w10892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10884w10896w10897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10889w10901w10902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10750w10766w10767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10894w10906w10907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10899w10911w10912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10904w10914w10915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10909w10917w10918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10758w10771w10772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10764w10776w10777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10769w10781w10782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10774w10786w10787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10779w10791w10792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10784w10796w10797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10789w10801w10802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range458w461w462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range463w466w467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range468w471w472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range473w476w477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range478w481w482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range483w486w487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range488w491w492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range493w496w497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range498w501w502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range503w506w507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range508w511w512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range513w516w517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range518w521w522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range523w526w527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range528w531w532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range533w536w537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range538w541w542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range543w546w547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range548w551w552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range553w556w557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range418w421w422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range558w561w562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range563w566w567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range568w571w572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range573w576w577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range423w426w427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range428w431w432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range433w436w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range438w441w442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range443w446w447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range448w451w452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range453w456w457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7570w7784w7785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7629w7866w7867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7635w7874w7875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7641w7882w7883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7647w7890w7891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7653w7898w7899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7659w7906w7907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7665w7914w7915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7671w7922w7923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7677w7930w7931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7683w7938w7939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7575w7794w7795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7689w7946w7947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7695w7954w7955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7701w7962w7963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7707w7970w7971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7711w7978w7979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7523w7986w7987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7528w7994w7995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7530w8002w8003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7532w8010w8011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7534w8018w8019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7581w7802w7803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7536w8026w8027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7538w8034w8035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7540w8042w8043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7542w8050w8051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7587w7810w7811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7593w7818w7819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7599w7826w7827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7605w7834w7835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7611w7842w7843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7617w7850w7851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7623w7858w7859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8386w8591w8592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8445w8673w8674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8451w8681w8682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8457w8689w8690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8463w8697w8698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8469w8705w8706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8475w8713w8714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8481w8721w8722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8487w8729w8730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8493w8737w8738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8499w8745w8746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8391w8601w8602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8505w8753w8754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8511w8761w8762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8517w8769w8770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8521w8777w8778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8335w8785w8786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8340w8793w8794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8342w8801w8802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8344w8809w8810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8346w8817w8818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8348w8825w8826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8397w8609w8610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8350w8833w8834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8352w8841w8842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8354w8849w8850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8356w8857w8858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8403w8617w8618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8409w8625w8626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8415w8633w8634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8421w8641w8642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8427w8649w8650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8433w8657w8658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8439w8665w8666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9197w9393w9394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9256w9475w9476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9262w9483w9484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9268w9491w9492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9274w9499w9500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9280w9507w9508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9286w9515w9516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9292w9523w9524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9298w9531w9532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9304w9539w9540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9310w9547w9548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9202w9403w9404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9316w9555w9556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9322w9563w9564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9326w9571w9572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9142w9579w9580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9147w9587w9588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9149w9595w9596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9151w9603w9604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9153w9611w9612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9155w9619w9620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9157w9627w9628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9208w9411w9412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9159w9635w9636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9161w9643w9644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9163w9651w9652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9165w9659w9660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9214w9419w9420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9220w9427w9428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9226w9435w9436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9232w9443w9444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9238w9451w9452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9244w9459w9460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9250w9467w9468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range862w1148w1149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range921w1230w1231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range927w1238w1239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range933w1246w1247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range939w1254w1255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range945w1262w1263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range951w1270w1271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range957w1278w1279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range963w1286w1287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range969w1294w1295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range975w1302w1303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range867w1158w1159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range981w1310w1311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range987w1318w1319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range993w1326w1327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range999w1334w1335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1005w1342w1343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1011w1350w1351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1017w1358w1359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1023w1366w1367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1029w1374w1375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1035w1382w1383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range873w1166w1167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1041w1390w1391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1047w1398w1399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1051w1406w1407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range847w1414w1415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range879w1174w1175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range885w1182w1183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range891w1190w1191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range897w1198w1199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range903w1206w1207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range909w1214w1215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range915w1222w1223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1718w1995w1996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1777w2077w2078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1783w2085w2086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1789w2093w2094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1795w2101w2102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1801w2109w2110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1807w2117w2118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1813w2125w2126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1819w2133w2134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1825w2141w2142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1831w2149w2150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1723w2005w2006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1837w2157w2158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1843w2165w2166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1849w2173w2174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1855w2181w2182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1861w2189w2190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1867w2197w2198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1873w2205w2206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1879w2213w2214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1885w2221w2222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1891w2229w2230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1729w2013w2014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1897w2237w2238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1901w2245w2246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1699w2253w2254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1704w2261w2262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1735w2021w2022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1741w2029w2030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1747w2037w2038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1753w2045w2046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1759w2053w2054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1765w2061w2062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1771w2069w2070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2569w2837w2838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2628w2919w2920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2634w2927w2928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2640w2935w2936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2646w2943w2944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2652w2951w2952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2658w2959w2960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2664w2967w2968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2670w2975w2976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2676w2983w2984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2682w2991w2992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2574w2847w2848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2688w2999w3000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2694w3007w3008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2700w3015w3016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2706w3023w3024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2712w3031w3032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2718w3039w3040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2724w3047w3048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2730w3055w3056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2736w3063w3064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2742w3071w3072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2580w2855w2856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2746w3079w3080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2546w3087w3088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2551w3095w3096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2553w3103w3104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2586w2863w2864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2592w2871w2872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2598w2879w2880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2604w2887w2888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2610w2895w2896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2616w2903w2904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2622w2911w2912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3415w3674w3675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3474w3756w3757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3480w3764w3765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3486w3772w3773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3492w3780w3781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3498w3788w3789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3504w3796w3797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3510w3804w3805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3516w3812w3813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3522w3820w3821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3528w3828w3829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3420w3684w3685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3534w3836w3837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3540w3844w3845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3546w3852w3853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3552w3860w3861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3558w3868w3869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3564w3876w3877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3570w3884w3885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3576w3892w3893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3582w3900w3901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3586w3908w3909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3426w3692w3693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3388w3916w3917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3393w3924w3925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3395w3932w3933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3397w3940w3941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3432w3700w3701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3438w3708w3709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3444w3716w3717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3450w3724w3725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3456w3732w3733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3462w3740w3741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3468w3748w3749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4256w4506w4507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4315w4588w4589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4321w4596w4597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4327w4604w4605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4333w4612w4613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4339w4620w4621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4345w4628w4629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4351w4636w4637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4357w4644w4645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4363w4652w4653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4369w4660w4661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4261w4516w4517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4375w4668w4669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4381w4676w4677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4387w4684w4685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4393w4692w4693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4399w4700w4701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4405w4708w4709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4411w4716w4717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4417w4724w4725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4421w4732w4733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4225w4740w4741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4267w4524w4525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4230w4748w4749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4232w4756w4757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4234w4764w4765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4236w4772w4773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4273w4532w4533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4279w4540w4541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4285w4548w4549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4291w4556w4557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4297w4564w4565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4303w4572w4573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4309w4580w4581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5092w5333w5334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5151w5415w5416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5157w5423w5424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5163w5431w5432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5169w5439w5440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5175w5447w5448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5181w5455w5456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5187w5463w5464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5193w5471w5472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5199w5479w5480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5205w5487w5488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5097w5343w5344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5211w5495w5496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5217w5503w5504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5223w5511w5512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5229w5519w5520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5235w5527w5528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5241w5535w5536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5247w5543w5544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5251w5551w5552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5057w5559w5560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5062w5567w5568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5103w5351w5352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5064w5575w5576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5066w5583w5584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5068w5591w5592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5070w5599w5600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5109w5359w5360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5115w5367w5368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5121w5375w5376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5127w5383w5384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5133w5391w5392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5139w5399w5400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5145w5407w5408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5923w6155w6156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5982w6237w6238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5988w6245w6246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5994w6253w6254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6000w6261w6262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6006w6269w6270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6012w6277w6278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6018w6285w6286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6024w6293w6294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6030w6301w6302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6036w6309w6310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5928w6165w6166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6042w6317w6318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6048w6325w6326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6054w6333w6334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6060w6341w6342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6066w6349w6350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6072w6357w6358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6076w6365w6366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5884w6373w6374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5889w6381w6382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5891w6389w6390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5934w6173w6174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5893w6397w6398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5895w6405w6406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5897w6413w6414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5899w6421w6422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5940w6181w6182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5946w6189w6190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5952w6197w6198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5958w6205w6206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5964w6213w6214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5970w6221w6222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5976w6229w6230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6749w6972w6973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6808w7054w7055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6814w7062w7063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6820w7070w7071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6826w7078w7079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6832w7086w7087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6838w7094w7095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6844w7102w7103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6850w7110w7111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6856w7118w7119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6862w7126w7127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6754w6982w6983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6868w7134w7135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6874w7142w7143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6880w7150w7151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6886w7158w7159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6892w7166w7167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6896w7174w7175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6706w7182w7183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6711w7190w7191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6713w7198w7199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6715w7206w7207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6760w6990w6991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6717w7214w7215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6719w7222w7223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6721w7230w7231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6723w7238w7239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6766w6998w6999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6772w7006w7007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6778w7014w7015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6784w7022w7023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6790w7030w7031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6796w7038w7039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6802w7046w7047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7572w7789w7790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7631w7870w7871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7637w7878w7879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7643w7886w7887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7649w7894w7895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7655w7902w7903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7661w7910w7911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7667w7918w7919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7673w7926w7927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7679w7934w7935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7685w7942w7943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7577w7798w7799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7691w7950w7951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7697w7958w7959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7703w7966w7967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7709w7974w7975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7712w7982w7983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7526w7990w7991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7529w7998w7999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7531w8006w8007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7533w8014w8015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7535w8022w8023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7583w7806w7807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7537w8030w8031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7539w8038w8039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7541w8046w8047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7543w8054w8055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7589w7814w7815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7595w7822w7823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7601w7830w7831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7607w7838w7839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7613w7846w7847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7619w7854w7855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7625w7862w7863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8388w8596w8597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8447w8677w8678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8453w8685w8686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8459w8693w8694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8465w8701w8702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8471w8709w8710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8477w8717w8718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8483w8725w8726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8489w8733w8734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8495w8741w8742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8501w8749w8750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8393w8605w8606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8507w8757w8758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8513w8765w8766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8519w8773w8774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8522w8781w8782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8338w8789w8790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8341w8797w8798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8343w8805w8806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8345w8813w8814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8347w8821w8822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8349w8829w8830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8399w8613w8614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8351w8837w8838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8353w8845w8846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8355w8853w8854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8357w8861w8862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8405w8621w8622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8411w8629w8630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8417w8637w8638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8423w8645w8646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8429w8653w8654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8435w8661w8662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8441w8669w8670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9199w9398w9399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9258w9479w9480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9264w9487w9488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9270w9495w9496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9276w9503w9504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9282w9511w9512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9288w9519w9520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9294w9527w9528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9300w9535w9536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9306w9543w9544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9312w9551w9552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9204w9407w9408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9318w9559w9560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9324w9567w9568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9327w9575w9576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9145w9583w9584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9148w9591w9592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9150w9599w9600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9152w9607w9608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9154w9615w9616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9156w9623w9624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9158w9631w9632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9210w9415w9416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9160w9639w9640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9162w9647w9648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9164w9655w9656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9166w9663w9664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9216w9423w9424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9222w9431w9432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9228w9439w9440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9234w9447w9448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9240w9455w9456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9246w9463w9464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9252w9471w9472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w10269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range864w1153w1154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range923w1234w1235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range929w1242w1243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range935w1250w1251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range941w1258w1259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range947w1266w1267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range953w1274w1275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range959w1282w1283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range965w1290w1291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range971w1298w1299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range977w1306w1307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range869w1162w1163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range983w1314w1315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range989w1322w1323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range995w1330w1331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1001w1338w1339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1007w1346w1347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1013w1354w1355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1019w1362w1363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1025w1370w1371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1031w1378w1379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1037w1386w1387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range875w1170w1171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1043w1394w1395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1049w1402w1403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1052w1410w1411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range850w1418w1419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range881w1178w1179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range887w1186w1187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range893w1194w1195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range899w1202w1203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range905w1210w1211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range911w1218w1219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range917w1226w1227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1720w2000w2001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1779w2081w2082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1785w2089w2090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1791w2097w2098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1797w2105w2106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1803w2113w2114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1809w2121w2122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1815w2129w2130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1821w2137w2138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1827w2145w2146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1833w2153w2154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1725w2009w2010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1839w2161w2162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1845w2169w2170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1851w2177w2178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1857w2185w2186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1863w2193w2194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1869w2201w2202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1875w2209w2210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1881w2217w2218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1887w2225w2226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1893w2233w2234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1731w2017w2018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1899w2241w2242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1902w2249w2250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1702w2257w2258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1705w2265w2266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1737w2025w2026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1743w2033w2034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1749w2041w2042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1755w2049w2050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1761w2057w2058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1767w2065w2066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1773w2073w2074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2571w2842w2843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2630w2923w2924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2636w2931w2932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2642w2939w2940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2648w2947w2948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2654w2955w2956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2660w2963w2964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2666w2971w2972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2672w2979w2980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2678w2987w2988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2684w2995w2996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2576w2851w2852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2690w3003w3004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2696w3011w3012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2702w3019w3020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2708w3027w3028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2714w3035w3036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2720w3043w3044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2726w3051w3052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2732w3059w3060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2738w3067w3068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2744w3075w3076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2582w2859w2860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2747w3083w3084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2549w3091w3092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2552w3099w3100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2554w3107w3108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2588w2867w2868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2594w2875w2876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2600w2883w2884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2606w2891w2892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2612w2899w2900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2618w2907w2908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2624w2915w2916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3417w3679w3680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3476w3760w3761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3482w3768w3769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3488w3776w3777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3494w3784w3785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3500w3792w3793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3506w3800w3801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3512w3808w3809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3518w3816w3817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3524w3824w3825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3530w3832w3833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3422w3688w3689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3536w3840w3841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3542w3848w3849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3548w3856w3857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3554w3864w3865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3560w3872w3873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3566w3880w3881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3572w3888w3889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3578w3896w3897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3584w3904w3905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3587w3912w3913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3428w3696w3697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3391w3920w3921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3394w3928w3929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3396w3936w3937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3398w3944w3945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3434w3704w3705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3440w3712w3713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3446w3720w3721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3452w3728w3729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3458w3736w3737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3464w3744w3745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3470w3752w3753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4258w4511w4512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4317w4592w4593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4323w4600w4601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4329w4608w4609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4335w4616w4617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4341w4624w4625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4347w4632w4633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4353w4640w4641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4359w4648w4649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4365w4656w4657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4371w4664w4665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4263w4520w4521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4377w4672w4673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4383w4680w4681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4389w4688w4689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4395w4696w4697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4401w4704w4705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4407w4712w4713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4413w4720w4721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4419w4728w4729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4422w4736w4737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4228w4744w4745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4269w4528w4529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4231w4752w4753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4233w4760w4761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4235w4768w4769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4237w4776w4777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4275w4536w4537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4281w4544w4545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4287w4552w4553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4293w4560w4561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4299w4568w4569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4305w4576w4577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4311w4584w4585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5094w5338w5339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5153w5419w5420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5159w5427w5428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5165w5435w5436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5171w5443w5444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5177w5451w5452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5183w5459w5460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5189w5467w5468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5195w5475w5476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5201w5483w5484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5207w5491w5492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5099w5347w5348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5213w5499w5500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5219w5507w5508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5225w5515w5516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5231w5523w5524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5237w5531w5532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5243w5539w5540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5249w5547w5548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5252w5555w5556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5060w5563w5564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5063w5571w5572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5105w5355w5356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5065w5579w5580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5067w5587w5588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5069w5595w5596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5071w5603w5604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5111w5363w5364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5117w5371w5372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5123w5379w5380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5129w5387w5388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5135w5395w5396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5141w5403w5404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5147w5411w5412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5925w6160w6161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5984w6241w6242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5990w6249w6250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5996w6257w6258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6002w6265w6266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6008w6273w6274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6014w6281w6282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6020w6289w6290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6026w6297w6298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6032w6305w6306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6038w6313w6314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5930w6169w6170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6044w6321w6322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6050w6329w6330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6056w6337w6338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6062w6345w6346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6068w6353w6354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6074w6361w6362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6077w6369w6370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5887w6377w6378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5890w6385w6386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5892w6393w6394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5936w6177w6178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5894w6401w6402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5896w6409w6410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5898w6417w6418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5900w6425w6426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5942w6185w6186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5948w6193w6194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5954w6201w6202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5960w6209w6210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5966w6217w6218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5972w6225w6226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5978w6233w6234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6751w6977w6978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6810w7058w7059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6816w7066w7067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6822w7074w7075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6828w7082w7083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6834w7090w7091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6840w7098w7099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6846w7106w7107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6852w7114w7115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6858w7122w7123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6864w7130w7131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6756w6986w6987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6870w7138w7139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6876w7146w7147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6882w7154w7155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6888w7162w7163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6894w7170w7171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6897w7178w7179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6709w7186w7187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6712w7194w7195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6714w7202w7203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6716w7210w7211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6762w6994w6995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6718w7218w7219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6720w7226w7227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6722w7234w7235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6724w7242w7243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6768w7002w7003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6774w7010w7011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6780w7018w7019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6786w7026w7027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6792w7034w7035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6798w7042w7043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6804w7050w7051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8871w8872w8873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8952w8953w8954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8960w8961w8962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8968w8969w8970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8976w8977w8978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8984w8985w8986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8992w8993w8994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9000w9001w9002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9008w9009w9010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9016w9017w9018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9024w9025w9026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8880w8881w8882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9032w9033w9034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9040w9041w9042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9048w9049w9050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9056w9057w9058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9064w9065w9066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9072w9073w9074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9080w9081w9082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9088w9089w9090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9096w9097w9098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9104w9105w9106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8888w8889w8890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9112w9113w9114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9120w9121w9122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9128w9129w9130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9136w9137w9138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8896w8897w8898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8904w8905w8906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8912w8913w8914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8920w8921w8922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8928w8929w8930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8936w8937w8938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8944w8945w8946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9673w9674w9675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9754w9755w9756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9762w9763w9764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9770w9771w9772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9778w9779w9780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9786w9787w9788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9794w9795w9796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9802w9803w9804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9810w9811w9812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9818w9819w9820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9826w9827w9828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9682w9683w9684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9834w9835w9836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9842w9843w9844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9850w9851w9852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9858w9859w9860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9866w9867w9868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9874w9875w9876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9882w9883w9884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9890w9891w9892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9898w9899w9900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9906w9907w9908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9690w9691w9692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9914w9915w9916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9922w9923w9924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9930w9931w9932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9938w9939w9940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9698w9699w9700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9706w9707w9708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9714w9715w9716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9722w9723w9724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9730w9731w9732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9738w9739w9740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9746w9747w9748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10470w10471w10472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10551w10552w10553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10559w10560w10561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10567w10568w10569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10575w10576w10577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10583w10584w10585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10591w10592w10593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10599w10600w10601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10607w10608w10609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10615w10616w10617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10623w10624w10625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10479w10480w10481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10631w10632w10633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10639w10640w10641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10647w10648w10649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10655w10656w10657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10663w10664w10665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10671w10672w10673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10679w10680w10681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10687w10688w10689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10695w10696w10697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10703w10704w10705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10487w10488w10489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10711w10712w10713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10719w10720w10721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10727w10728w10729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10735w10736w10737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10495w10496w10497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10503w10504w10505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10511w10512w10513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10519w10520w10521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10527w10528w10529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10535w10536w10537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10543w10544w10545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1428w1429w1430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1509w1510w1511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1517w1518w1519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1525w1526w1527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1533w1534w1535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1541w1542w1543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1549w1550w1551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1557w1558w1559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1565w1566w1567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1573w1574w1575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1581w1582w1583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1437w1438w1439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1589w1590w1591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1597w1598w1599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1605w1606w1607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1613w1614w1615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1621w1622w1623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1629w1630w1631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1637w1638w1639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1645w1646w1647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1653w1654w1655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1661w1662w1663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1445w1446w1447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1669w1670w1671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1677w1678w1679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1685w1686w1687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1693w1694w1695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1453w1454w1455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1461w1462w1463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1469w1470w1471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1477w1478w1479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1485w1486w1487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1493w1494w1495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1501w1502w1503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2275w2276w2277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2356w2357w2358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2364w2365w2366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2372w2373w2374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2380w2381w2382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2388w2389w2390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2396w2397w2398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2404w2405w2406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2412w2413w2414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2420w2421w2422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2428w2429w2430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2284w2285w2286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2436w2437w2438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2444w2445w2446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2452w2453w2454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2460w2461w2462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2468w2469w2470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2476w2477w2478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2484w2485w2486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2492w2493w2494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2500w2501w2502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2508w2509w2510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2292w2293w2294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2516w2517w2518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2524w2525w2526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2532w2533w2534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2540w2541w2542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2300w2301w2302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2308w2309w2310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2316w2317w2318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2324w2325w2326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2332w2333w2334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2340w2341w2342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2348w2349w2350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3117w3118w3119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3198w3199w3200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3206w3207w3208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3214w3215w3216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3222w3223w3224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3230w3231w3232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3238w3239w3240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3246w3247w3248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3254w3255w3256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3262w3263w3264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3270w3271w3272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3126w3127w3128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3278w3279w3280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3286w3287w3288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3294w3295w3296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3302w3303w3304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3310w3311w3312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3318w3319w3320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3326w3327w3328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3334w3335w3336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3342w3343w3344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3350w3351w3352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3134w3135w3136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3358w3359w3360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3366w3367w3368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3374w3375w3376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3382w3383w3384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3142w3143w3144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3150w3151w3152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3158w3159w3160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3166w3167w3168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3174w3175w3176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3182w3183w3184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3190w3191w3192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3954w3955w3956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4035w4036w4037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4043w4044w4045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4051w4052w4053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4059w4060w4061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4067w4068w4069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4075w4076w4077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4083w4084w4085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4091w4092w4093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4099w4100w4101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4107w4108w4109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3963w3964w3965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4115w4116w4117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4123w4124w4125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4131w4132w4133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4139w4140w4141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4147w4148w4149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4155w4156w4157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4163w4164w4165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4171w4172w4173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4179w4180w4181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4187w4188w4189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3971w3972w3973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4195w4196w4197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4203w4204w4205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4211w4212w4213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4219w4220w4221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3979w3980w3981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3987w3988w3989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3995w3996w3997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4003w4004w4005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4011w4012w4013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4019w4020w4021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4027w4028w4029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4786w4787w4788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4867w4868w4869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4875w4876w4877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4883w4884w4885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4891w4892w4893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4899w4900w4901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4907w4908w4909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4915w4916w4917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4923w4924w4925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4931w4932w4933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4939w4940w4941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4795w4796w4797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4947w4948w4949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4955w4956w4957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4963w4964w4965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4971w4972w4973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4979w4980w4981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4987w4988w4989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4995w4996w4997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5003w5004w5005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5011w5012w5013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5019w5020w5021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4803w4804w4805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5027w5028w5029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5035w5036w5037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5043w5044w5045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5051w5052w5053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4811w4812w4813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4819w4820w4821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4827w4828w4829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4835w4836w4837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4843w4844w4845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4851w4852w4853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4859w4860w4861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5613w5614w5615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5694w5695w5696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5702w5703w5704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5710w5711w5712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5718w5719w5720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5726w5727w5728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5734w5735w5736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5742w5743w5744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5750w5751w5752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5758w5759w5760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5766w5767w5768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5622w5623w5624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5774w5775w5776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5782w5783w5784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5790w5791w5792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5798w5799w5800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5806w5807w5808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5814w5815w5816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5822w5823w5824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5830w5831w5832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5838w5839w5840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5846w5847w5848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5630w5631w5632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5854w5855w5856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5862w5863w5864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5870w5871w5872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5878w5879w5880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5638w5639w5640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5646w5647w5648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5654w5655w5656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5662w5663w5664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5670w5671w5672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5678w5679w5680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5686w5687w5688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6435w6436w6437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6516w6517w6518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6524w6525w6526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6532w6533w6534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6540w6541w6542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6548w6549w6550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6556w6557w6558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6564w6565w6566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6572w6573w6574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6580w6581w6582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6588w6589w6590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6444w6445w6446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6596w6597w6598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6604w6605w6606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6612w6613w6614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6620w6621w6622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6628w6629w6630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6636w6637w6638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6644w6645w6646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6652w6653w6654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6660w6661w6662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6668w6669w6670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6452w6453w6454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6676w6677w6678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6684w6685w6686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6692w6693w6694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6700w6701w6702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6460w6461w6462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6468w6469w6470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6476w6477w6478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6484w6485w6486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6492w6493w6494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6500w6501w6502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6508w6509w6510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7252w7253w7254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7333w7334w7335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7341w7342w7343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7349w7350w7351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7357w7358w7359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7365w7366w7367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7373w7374w7375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7381w7382w7383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7389w7390w7391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7397w7398w7399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7405w7406w7407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7261w7262w7263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7413w7414w7415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7421w7422w7423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7429w7430w7431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7437w7438w7439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7445w7446w7447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7453w7454w7455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7461w7462w7463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7469w7470w7471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7477w7478w7479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7485w7486w7487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7269w7270w7271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7493w7494w7495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7501w7502w7503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7509w7510w7511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7517w7518w7519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7277w7278w7279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7285w7286w7287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7293w7294w7295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7301w7302w7303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7309w7310w7311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7317w7318w7319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7325w7326w7327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8064w8065w8066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8145w8146w8147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8153w8154w8155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8161w8162w8163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8169w8170w8171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8177w8178w8179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8185w8186w8187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8193w8194w8195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8201w8202w8203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8209w8210w8211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8217w8218w8219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8073w8074w8075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8225w8226w8227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8233w8234w8235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8241w8242w8243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8249w8250w8251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8257w8258w8259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8265w8266w8267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8273w8274w8275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8281w8282w8283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8289w8290w8291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8297w8298w8299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8081w8082w8083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8305w8306w8307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8313w8314w8315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8321w8322w8323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8329w8330w8331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8089w8090w8091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8097w8098w8099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8105w8106w8107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8113w8114w8115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8121w8122w8123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8129w8130w8131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8137w8138w8139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_estimate_w10920w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7786w8058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7868w8141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7876w8149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7884w8157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7892w8165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7900w8173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7908w8181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7916w8189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7924w8197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7932w8205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7940w8213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7796w8069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7948w8221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7956w8229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7964w8237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7972w8245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7980w8253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7988w8261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7996w8269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8004w8277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8012w8285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8020w8293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7804w8077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8028w8301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8036w8309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8044w8317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8052w8325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7812w8085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7820w8093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7828w8101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7836w8109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7844w8117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7852w8125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7860w8133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8593w8865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8675w8948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8683w8956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8691w8964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8699w8972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8707w8980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8715w8988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8723w8996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8731w9004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8739w9012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8747w9020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8603w8876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8755w9028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8763w9036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8771w9044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8779w9052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8787w9060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8795w9068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8803w9076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8811w9084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8819w9092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8827w9100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8611w8884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8835w9108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8843w9116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8851w9124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8859w9132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8619w8892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8627w8900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8635w8908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8643w8916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8651w8924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8659w8932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8667w8940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9395w9667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9477w9750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9485w9758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9493w9766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9501w9774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9509w9782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9517w9790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9525w9798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9533w9806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9541w9814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9549w9822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9405w9678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9557w9830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9565w9838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9573w9846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9581w9854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9589w9862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9597w9870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9605w9878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9613w9886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9621w9894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9629w9902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9413w9686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9637w9910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9645w9918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9653w9926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9661w9934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9421w9694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9429w9702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9437w9710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9445w9718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9453w9726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9461w9734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9469w9742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10192w10464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10274w10547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10282w10555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10290w10563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10298w10571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10306w10579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10314w10587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10322w10595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10330w10603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10338w10611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10346w10619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10202w10475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10354w10627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10362w10635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10370w10643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10378w10651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10386w10659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10394w10667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10402w10675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10410w10683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10418w10691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10426w10699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10210w10483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10434w10707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10442w10715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10450w10723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10458w10731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10218w10491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10226w10499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10234w10507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10242w10515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10250w10523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10258w10531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10266w10539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1150w1422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1232w1505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1240w1513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1248w1521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1256w1529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1264w1537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1272w1545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1280w1553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1288w1561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1296w1569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1304w1577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1160w1433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1312w1585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1320w1593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1328w1601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1336w1609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1344w1617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1352w1625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1360w1633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1368w1641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1376w1649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1384w1657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1168w1441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1392w1665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1400w1673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1408w1681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1416w1689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1176w1449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1184w1457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1192w1465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1200w1473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1208w1481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1216w1489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1224w1497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1997w2269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2079w2352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2087w2360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2095w2368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2103w2376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2111w2384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2119w2392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2127w2400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2135w2408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2143w2416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2151w2424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2007w2280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2159w2432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2167w2440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2175w2448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2183w2456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2191w2464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2199w2472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2207w2480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2215w2488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2223w2496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2231w2504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2015w2288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2239w2512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2247w2520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2255w2528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2263w2536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2023w2296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2031w2304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2039w2312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2047w2320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2055w2328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2063w2336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2071w2344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2839w3111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2921w3194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2929w3202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2937w3210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2945w3218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2953w3226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2961w3234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2969w3242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2977w3250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2985w3258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2993w3266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2849w3122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3001w3274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3009w3282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3017w3290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3025w3298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3033w3306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3041w3314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3049w3322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3057w3330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3065w3338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3073w3346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2857w3130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3081w3354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3089w3362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3097w3370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3105w3378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2865w3138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2873w3146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2881w3154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2889w3162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2897w3170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2905w3178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2913w3186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3676w3948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3758w4031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3766w4039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3774w4047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3782w4055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3790w4063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3798w4071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3806w4079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3814w4087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3822w4095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3830w4103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3686w3959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3838w4111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3846w4119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3854w4127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3862w4135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3870w4143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3878w4151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3886w4159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3894w4167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3902w4175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3910w4183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3694w3967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3918w4191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3926w4199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3934w4207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3942w4215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3702w3975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3710w3983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3718w3991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3726w3999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3734w4007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3742w4015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3750w4023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4508w4780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4590w4863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4598w4871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4606w4879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4614w4887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4622w4895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4630w4903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4638w4911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4646w4919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4654w4927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4662w4935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4518w4791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4670w4943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4678w4951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4686w4959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4694w4967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4702w4975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4710w4983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4718w4991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4726w4999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4734w5007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4742w5015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4526w4799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4750w5023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4758w5031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4766w5039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4774w5047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4534w4807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4542w4815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4550w4823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4558w4831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4566w4839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4574w4847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4582w4855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5335w5607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5417w5690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5425w5698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5433w5706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5441w5714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5449w5722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5457w5730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5465w5738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5473w5746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5481w5754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5489w5762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5345w5618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5497w5770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5505w5778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5513w5786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5521w5794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5529w5802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5537w5810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5545w5818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5553w5826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5561w5834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5569w5842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5353w5626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5577w5850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5585w5858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5593w5866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5601w5874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5361w5634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5369w5642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5377w5650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5385w5658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5393w5666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5401w5674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5409w5682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6157w6429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6239w6512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6247w6520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6255w6528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6263w6536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6271w6544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6279w6552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6287w6560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6295w6568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6303w6576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6311w6584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6167w6440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6319w6592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6327w6600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6335w6608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6343w6616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6351w6624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6359w6632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6367w6640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6375w6648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6383w6656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6391w6664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6175w6448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6399w6672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6407w6680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6415w6688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6423w6696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6183w6456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6191w6464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6199w6472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6207w6480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6215w6488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6223w6496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6231w6504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6974w7246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7056w7329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7064w7337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7072w7345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7080w7353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7088w7361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7096w7369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7104w7377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7112w7385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7120w7393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7128w7401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6984w7257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7136w7409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7144w7417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7152w7425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7160w7433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7168w7441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7176w7449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7184w7457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7192w7465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7200w7473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7208w7481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6992w7265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7216w7489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7224w7497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7232w7505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7240w7513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7000w7273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7008w7281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7016w7289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7024w7297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7032w7305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7040w7313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7048w7321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7791w8061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7872w8143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7880w8151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7888w8159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7896w8167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7904w8175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7912w8183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7920w8191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7928w8199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7936w8207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7944w8215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7800w8071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7952w8223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7960w8231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7968w8239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7976w8247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7984w8255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7992w8263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8000w8271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8008w8279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8016w8287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8024w8295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7808w8079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8032w8303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8040w8311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8048w8319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8056w8327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7816w8087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7824w8095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7832w8103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7840w8111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7848w8119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7856w8127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7864w8135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8598w8868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8679w8950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8687w8958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8695w8966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8703w8974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8711w8982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8719w8990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8727w8998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8735w9006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8743w9014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8751w9022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8607w8878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8759w9030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8767w9038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8775w9046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8783w9054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8791w9062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8799w9070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8807w9078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8815w9086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8823w9094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8831w9102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8615w8886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8839w9110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8847w9118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8855w9126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8863w9134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8623w8894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8631w8902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8639w8910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8647w8918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8655w8926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8663w8934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8671w8942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9400w9670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9481w9752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9489w9760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9497w9768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9505w9776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9513w9784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9521w9792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9529w9800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9537w9808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9545w9816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9553w9824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9409w9680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9561w9832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9569w9840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9577w9848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9585w9856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9593w9864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9601w9872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9609w9880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9617w9888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9625w9896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9633w9904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9417w9688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9641w9912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9649w9920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9657w9928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9665w9936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9425w9696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9433w9704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9441w9712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9449w9720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9457w9728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9465w9736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9473w9744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10197w10467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10278w10549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10286w10557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10294w10565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10302w10573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10310w10581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10318w10589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10326w10597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10334w10605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10342w10613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10350w10621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10206w10477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10358w10629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10366w10637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10374w10645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10382w10653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10390w10661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10398w10669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10406w10677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10414w10685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10422w10693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10430w10701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10214w10485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10438w10709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10446w10717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10454w10725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10462w10733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10222w10493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10230w10501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10238w10509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10246w10517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10254w10525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10262w10533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10270w10541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1155w1425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1236w1507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1244w1515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1252w1523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1260w1531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1268w1539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1276w1547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1284w1555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1292w1563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1300w1571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1308w1579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1164w1435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1316w1587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1324w1595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1332w1603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1340w1611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1348w1619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1356w1627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1364w1635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1372w1643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1380w1651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1388w1659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1172w1443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1396w1667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1404w1675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1412w1683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1420w1691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1180w1451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1188w1459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1196w1467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1204w1475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1212w1483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1220w1491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1228w1499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2002w2272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2083w2354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2091w2362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2099w2370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2107w2378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2115w2386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2123w2394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2131w2402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2139w2410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2147w2418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2155w2426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2011w2282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2163w2434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2171w2442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2179w2450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2187w2458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2195w2466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2203w2474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2211w2482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2219w2490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2227w2498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2235w2506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2019w2290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2243w2514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2251w2522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2259w2530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2267w2538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2027w2298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2035w2306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2043w2314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2051w2322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2059w2330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2067w2338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2075w2346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2844w3114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2925w3196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2933w3204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2941w3212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2949w3220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2957w3228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2965w3236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2973w3244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2981w3252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2989w3260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2997w3268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2853w3124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3005w3276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3013w3284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3021w3292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3029w3300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3037w3308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3045w3316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3053w3324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3061w3332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3069w3340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3077w3348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2861w3132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3085w3356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3093w3364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3101w3372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3109w3380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2869w3140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2877w3148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2885w3156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2893w3164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2901w3172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2909w3180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2917w3188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3681w3951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3762w4033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3770w4041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3778w4049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3786w4057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3794w4065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3802w4073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3810w4081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3818w4089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3826w4097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3834w4105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3690w3961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3842w4113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3850w4121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3858w4129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3866w4137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3874w4145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3882w4153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3890w4161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3898w4169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3906w4177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3914w4185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3698w3969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3922w4193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3930w4201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3938w4209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3946w4217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3706w3977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3714w3985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3722w3993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3730w4001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3738w4009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3746w4017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3754w4025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4513w4783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4594w4865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4602w4873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4610w4881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4618w4889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4626w4897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4634w4905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4642w4913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4650w4921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4658w4929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4666w4937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4522w4793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4674w4945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4682w4953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4690w4961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4698w4969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4706w4977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4714w4985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4722w4993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4730w5001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4738w5009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4746w5017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4530w4801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4754w5025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4762w5033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4770w5041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4778w5049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4538w4809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4546w4817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4554w4825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4562w4833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4570w4841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4578w4849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4586w4857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5340w5610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5421w5692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5429w5700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5437w5708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5445w5716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5453w5724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5461w5732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5469w5740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5477w5748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5485w5756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5493w5764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5349w5620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5501w5772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5509w5780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5517w5788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5525w5796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5533w5804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5541w5812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5549w5820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5557w5828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5565w5836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5573w5844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5357w5628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5581w5852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5589w5860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5597w5868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5605w5876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5365w5636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5373w5644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5381w5652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5389w5660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5397w5668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5405w5676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5413w5684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6162w6432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6243w6514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6251w6522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6259w6530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6267w6538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6275w6546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6283w6554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6291w6562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6299w6570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6307w6578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6315w6586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6171w6442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6323w6594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6331w6602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6339w6610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6347w6618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6355w6626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6363w6634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6371w6642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6379w6650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6387w6658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6395w6666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6179w6450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6403w6674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6411w6682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6419w6690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6427w6698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6187w6458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6195w6466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6203w6474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6211w6482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6219w6490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6227w6498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6235w6506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6979w7249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7060w7331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7068w7339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7076w7347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7084w7355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7092w7363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7100w7371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7108w7379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7116w7387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7124w7395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7132w7403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6988w7259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7140w7411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7148w7419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7156w7427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7164w7435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7172w7443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7180w7451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7188w7459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7196w7467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7204w7475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7212w7483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6996w7267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7220w7491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7228w7499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7236w7507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7244w7515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7004w7275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7012w7283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7020w7291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7028w7299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7036w7307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7044w7315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7052w7323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  atannode_0_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_1_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  atannode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  delay_input_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  delay_pipe_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  estimate_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  indexpointnum_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  multiplier_input_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  multipliernode_w :	STD_LOGIC_VECTOR (67 DOWNTO 0);
	 SIGNAL  post_estimate_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  pre_estimate_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  radians_load_node_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  startindex_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  x_pipenode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_pipenode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodeone_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_prenodetwo_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_start_node_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  x_subnode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_pipenode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodeone_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_prenodetwo_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_1_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  y_subnode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_pipenode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_10_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_11_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_12_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_13_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_2_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_3_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_4_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_5_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_6_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_7_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_8_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  z_subnode_9_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range9136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range10543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range4027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range5051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range7325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range8137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range8052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range9469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range10266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range3105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range6231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range7048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range8439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range9250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range10056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range1051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range5145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range6076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range8056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range9473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range10270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range3109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range6235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range7052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range8441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range9252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range10058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range1052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range5147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range6077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_45b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_l6b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_m6b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_n6b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_o6b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_55b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_65b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_75b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_85b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_95b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_a5b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_b5b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_c5b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_atan_d5b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_cordic_start_709
	 PORT
	 ( 
		index	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		value	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop30 : FOR i IN 0 TO 3 GENERATE 
		wire_ccc_cordic_m_w_lg_indexpointnum_w409w(i) <= indexpointnum_w(i) AND indexbit;
	END GENERATE loop30;
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10753w10754w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10753w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10794w10806w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10794w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10794w10795w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10794w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10799w10811w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10799w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10799w10800w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10799w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10804w10816w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10804w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10804w10805w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10804w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10809w10821w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10809w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10809w10810w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10809w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10814w10826w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10814w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10814w10815w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10814w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10819w10831w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10819w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10819w10820w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10819w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10824w10836w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10824w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10824w10825w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10824w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10829w10841w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10829w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10829w10830w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10829w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10834w10846w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10834w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10834w10835w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10834w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10839w10851w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10839w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10839w10840w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10839w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10760w10761w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10760w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10844w10856w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10844w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10844w10845w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10844w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10849w10861w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10849w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10849w10850w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10849w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10854w10866w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10854w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10854w10855w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10854w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10859w10871w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10859w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10859w10860w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10859w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10864w10876w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10864w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10864w10865w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10864w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10869w10881w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10869w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10869w10870w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10869w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10874w10886w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10874w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10874w10875w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10874w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10879w10891w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10879w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10879w10880w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10879w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10884w10896w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10884w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10884w10885w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10884w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10889w10901w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10889w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10889w10890w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10889w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10750w10766w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10750w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10750w10751w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10750w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10894w10906w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10894w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10894w10895w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10894w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10899w10911w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10899w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10899w10900w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10899w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10904w10914w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10904w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10904w10905w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10904w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10917w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10909w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10910w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10909w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10758w10771w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10758w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10758w10759w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10758w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10764w10776w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10764w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10764w10765w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10764w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10769w10781w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10769w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10769w10770w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10769w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10774w10786w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10774w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10774w10775w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10774w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10779w10791w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10779w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10779w10780w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10779w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10784w10796w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10784w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10784w10785w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10784w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10789w10801w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10789w(0) AND wire_indexbitff_w_lg_w_q_range10749w10752w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10789w10790w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10789w(0) AND wire_indexbitff_w_q_range10749w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range410w413w(0) <= wire_ccc_cordic_m_w_radians_range410w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range410w420w(0) <= wire_ccc_cordic_m_w_radians_range410w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range458w461w(0) <= wire_ccc_cordic_m_w_radians_range458w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range458w470w(0) <= wire_ccc_cordic_m_w_radians_range458w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range463w466w(0) <= wire_ccc_cordic_m_w_radians_range463w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range463w475w(0) <= wire_ccc_cordic_m_w_radians_range463w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range468w471w(0) <= wire_ccc_cordic_m_w_radians_range468w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range468w480w(0) <= wire_ccc_cordic_m_w_radians_range468w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range473w476w(0) <= wire_ccc_cordic_m_w_radians_range473w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range473w485w(0) <= wire_ccc_cordic_m_w_radians_range473w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range478w481w(0) <= wire_ccc_cordic_m_w_radians_range478w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range478w490w(0) <= wire_ccc_cordic_m_w_radians_range478w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range483w486w(0) <= wire_ccc_cordic_m_w_radians_range483w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range483w495w(0) <= wire_ccc_cordic_m_w_radians_range483w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range488w491w(0) <= wire_ccc_cordic_m_w_radians_range488w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range488w500w(0) <= wire_ccc_cordic_m_w_radians_range488w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range493w496w(0) <= wire_ccc_cordic_m_w_radians_range493w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range493w505w(0) <= wire_ccc_cordic_m_w_radians_range493w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range498w501w(0) <= wire_ccc_cordic_m_w_radians_range498w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range498w510w(0) <= wire_ccc_cordic_m_w_radians_range498w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range503w506w(0) <= wire_ccc_cordic_m_w_radians_range503w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range503w515w(0) <= wire_ccc_cordic_m_w_radians_range503w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range415w417w(0) <= wire_ccc_cordic_m_w_radians_range415w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range415w425w(0) <= wire_ccc_cordic_m_w_radians_range415w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range508w511w(0) <= wire_ccc_cordic_m_w_radians_range508w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range508w520w(0) <= wire_ccc_cordic_m_w_radians_range508w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range513w516w(0) <= wire_ccc_cordic_m_w_radians_range513w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range513w525w(0) <= wire_ccc_cordic_m_w_radians_range513w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range518w521w(0) <= wire_ccc_cordic_m_w_radians_range518w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range518w530w(0) <= wire_ccc_cordic_m_w_radians_range518w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range523w526w(0) <= wire_ccc_cordic_m_w_radians_range523w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range523w535w(0) <= wire_ccc_cordic_m_w_radians_range523w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range528w531w(0) <= wire_ccc_cordic_m_w_radians_range528w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range528w540w(0) <= wire_ccc_cordic_m_w_radians_range528w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range533w536w(0) <= wire_ccc_cordic_m_w_radians_range533w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range533w545w(0) <= wire_ccc_cordic_m_w_radians_range533w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range538w541w(0) <= wire_ccc_cordic_m_w_radians_range538w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range538w550w(0) <= wire_ccc_cordic_m_w_radians_range538w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range543w546w(0) <= wire_ccc_cordic_m_w_radians_range543w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range543w555w(0) <= wire_ccc_cordic_m_w_radians_range543w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range548w551w(0) <= wire_ccc_cordic_m_w_radians_range548w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range548w560w(0) <= wire_ccc_cordic_m_w_radians_range548w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range553w556w(0) <= wire_ccc_cordic_m_w_radians_range553w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range553w565w(0) <= wire_ccc_cordic_m_w_radians_range553w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range418w421w(0) <= wire_ccc_cordic_m_w_radians_range418w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range418w430w(0) <= wire_ccc_cordic_m_w_radians_range418w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range558w561w(0) <= wire_ccc_cordic_m_w_radians_range558w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range558w570w(0) <= wire_ccc_cordic_m_w_radians_range558w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range563w566w(0) <= wire_ccc_cordic_m_w_radians_range563w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range563w575w(0) <= wire_ccc_cordic_m_w_radians_range563w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range568w571w(0) <= wire_ccc_cordic_m_w_radians_range568w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range573w576w(0) <= wire_ccc_cordic_m_w_radians_range573w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range423w426w(0) <= wire_ccc_cordic_m_w_radians_range423w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range423w435w(0) <= wire_ccc_cordic_m_w_radians_range423w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range428w431w(0) <= wire_ccc_cordic_m_w_radians_range428w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range428w440w(0) <= wire_ccc_cordic_m_w_radians_range428w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range433w436w(0) <= wire_ccc_cordic_m_w_radians_range433w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range433w445w(0) <= wire_ccc_cordic_m_w_radians_range433w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range438w441w(0) <= wire_ccc_cordic_m_w_radians_range438w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range438w450w(0) <= wire_ccc_cordic_m_w_radians_range438w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range443w446w(0) <= wire_ccc_cordic_m_w_radians_range443w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range443w455w(0) <= wire_ccc_cordic_m_w_radians_range443w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range448w451w(0) <= wire_ccc_cordic_m_w_radians_range448w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range448w460w(0) <= wire_ccc_cordic_m_w_radians_range448w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range453w456w(0) <= wire_ccc_cordic_m_w_radians_range453w(0) AND wire_ccc_cordic_m_w_lg_indexbit412w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range453w465w(0) <= wire_ccc_cordic_m_w_radians_range453w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7570w7784w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7570w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7629w7866w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7629w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7635w7874w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7635w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7641w7882w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7641w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7647w7890w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7647w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7653w7898w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7653w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7659w7906w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7659w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7665w7914w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7665w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7671w7922w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7671w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7677w7930w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7677w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7683w7938w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7683w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7575w7794w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7575w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7689w7946w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7689w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7695w7954w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7695w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7701w7962w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7701w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7707w7970w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7707w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7711w7978w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7711w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7523w7986w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7523w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7528w7994w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7528w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7530w8002w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7530w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7532w8010w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7532w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7534w8018w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7534w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7581w7802w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7581w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7536w8026w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7536w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7538w8034w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7538w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7540w8042w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7540w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7542w8050w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7542w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7587w7810w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7587w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7593w7818w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7593w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7599w7826w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7599w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7605w7834w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7605w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7611w7842w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7611w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7617w7850w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7617w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7623w7858w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7623w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8386w8591w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8386w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8445w8673w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8445w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8451w8681w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8451w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8457w8689w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8457w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8463w8697w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8463w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8469w8705w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8469w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8475w8713w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8475w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8481w8721w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8481w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8487w8729w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8487w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8493w8737w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8493w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8499w8745w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8499w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8391w8601w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8391w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8505w8753w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8505w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8511w8761w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8511w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8517w8769w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8517w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8521w8777w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8521w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8335w8785w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8335w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8340w8793w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8340w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8342w8801w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8342w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8344w8809w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8344w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8346w8817w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8346w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8348w8825w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8348w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8397w8609w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8397w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8350w8833w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8350w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8352w8841w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8352w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8354w8849w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8354w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8356w8857w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8356w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8403w8617w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8403w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8409w8625w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8409w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8415w8633w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8415w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8421w8641w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8421w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8427w8649w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8427w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8433w8657w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8433w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8439w8665w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range8439w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9197w9393w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9197w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9256w9475w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9256w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9262w9483w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9262w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9268w9491w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9268w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9274w9499w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9274w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9280w9507w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9280w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9286w9515w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9286w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9292w9523w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9292w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9298w9531w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9298w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9304w9539w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9304w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9310w9547w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9310w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9202w9403w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9202w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9316w9555w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9316w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9322w9563w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9322w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9326w9571w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9326w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9142w9579w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9142w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9147w9587w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9147w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9149w9595w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9149w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9151w9603w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9151w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9153w9611w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9153w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9155w9619w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9155w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9157w9627w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9157w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9208w9411w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9208w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9159w9635w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9159w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9161w9643w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9161w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9163w9651w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9163w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9165w9659w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9165w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9214w9419w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9214w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9220w9427w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9220w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9226w9435w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9226w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9232w9443w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9232w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9238w9451w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9238w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9244w9459w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9244w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9250w9467w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range9250w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10003w10190w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10003w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10062w10272w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10062w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10068w10280w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10068w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10074w10288w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10074w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10080w10296w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10080w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10086w10304w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10086w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10092w10312w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10092w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10098w10320w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10098w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10104w10328w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10104w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10110w10336w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10110w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10116w10344w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10116w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10008w10200w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10008w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10122w10352w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10122w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10126w10360w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10126w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9944w10368w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9944w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9949w10376w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9949w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9951w10384w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9951w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9953w10392w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9953w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9955w10400w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9955w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9957w10408w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9957w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9959w10416w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9959w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9961w10424w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9961w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10014w10208w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10014w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9963w10432w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9963w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9965w10440w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9965w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9967w10448w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9967w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9969w10456w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9969w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10020w10216w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10020w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10026w10224w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10026w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10032w10232w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10032w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10038w10240w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10038w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10044w10248w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10044w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10050w10256w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10050w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10056w10264w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range10056w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range862w1148w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range862w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range921w1230w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range921w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range927w1238w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range927w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range933w1246w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range933w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range939w1254w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range939w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range945w1262w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range945w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range951w1270w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range951w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range957w1278w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range957w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range963w1286w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range963w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range969w1294w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range969w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range975w1302w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range975w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range867w1158w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range867w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range981w1310w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range981w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range987w1318w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range987w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range993w1326w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range993w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range999w1334w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range999w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1005w1342w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1005w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1011w1350w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1011w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1017w1358w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1017w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1023w1366w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1023w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1029w1374w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1029w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1035w1382w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1035w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range873w1166w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range873w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1041w1390w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1041w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1047w1398w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1047w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1051w1406w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range1051w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range847w1414w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range847w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range879w1174w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range879w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range885w1182w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range885w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range891w1190w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range891w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range897w1198w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range897w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range903w1206w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range903w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range909w1214w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range909w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range915w1222w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range915w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1718w1995w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1718w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1777w2077w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1777w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1783w2085w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1783w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1789w2093w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1789w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1795w2101w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1795w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1801w2109w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1801w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1807w2117w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1807w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1813w2125w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1813w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1819w2133w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1819w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1825w2141w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1825w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1831w2149w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1831w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1723w2005w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1723w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1837w2157w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1837w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1843w2165w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1843w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1849w2173w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1849w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1855w2181w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1855w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1861w2189w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1861w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1867w2197w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1867w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1873w2205w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1873w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1879w2213w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1879w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1885w2221w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1885w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1891w2229w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1891w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1729w2013w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1729w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1897w2237w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1897w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1901w2245w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1901w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1699w2253w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1699w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1704w2261w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1704w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1735w2021w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1735w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1741w2029w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1741w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1747w2037w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1747w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1753w2045w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1753w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1759w2053w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1759w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1765w2061w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1765w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1771w2069w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1771w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2569w2837w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2569w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2628w2919w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2628w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2634w2927w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2634w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2640w2935w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2640w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2646w2943w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2646w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2652w2951w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2652w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2658w2959w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2658w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2664w2967w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2664w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2670w2975w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2670w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2676w2983w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2676w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2682w2991w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2682w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2574w2847w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2574w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2688w2999w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2688w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2694w3007w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2694w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2700w3015w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2700w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2706w3023w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2706w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2712w3031w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2712w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2718w3039w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2718w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2724w3047w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2724w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2730w3055w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2730w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2736w3063w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2736w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2742w3071w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2742w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2580w2855w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2580w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2746w3079w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2746w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2546w3087w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2546w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2551w3095w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2551w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2553w3103w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2553w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2586w2863w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2586w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2592w2871w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2592w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2598w2879w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2598w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2604w2887w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2604w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2610w2895w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2610w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2616w2903w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2616w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2622w2911w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2622w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3415w3674w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3415w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3474w3756w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3474w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3480w3764w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3480w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3486w3772w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3486w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3492w3780w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3492w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3498w3788w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3498w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3504w3796w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3504w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3510w3804w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3510w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3516w3812w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3516w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3522w3820w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3522w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3528w3828w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3528w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3420w3684w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3420w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3534w3836w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3534w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3540w3844w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3540w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3546w3852w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3546w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3552w3860w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3552w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3558w3868w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3558w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3564w3876w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3564w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3570w3884w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3570w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3576w3892w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3576w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3582w3900w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3582w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3586w3908w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3586w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3426w3692w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3426w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3388w3916w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3388w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3393w3924w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3393w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3395w3932w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3395w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3397w3940w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3397w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3432w3700w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3432w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3438w3708w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3438w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3444w3716w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3444w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3450w3724w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3450w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3456w3732w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3456w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3462w3740w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3462w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3468w3748w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3468w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4256w4506w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4256w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4315w4588w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4315w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4321w4596w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4321w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4327w4604w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4327w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4333w4612w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4333w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4339w4620w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4339w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4345w4628w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4345w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4351w4636w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4351w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4357w4644w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4357w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4363w4652w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4363w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4369w4660w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4369w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4261w4516w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4261w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4375w4668w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4375w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4381w4676w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4381w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4387w4684w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4387w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4393w4692w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4393w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4399w4700w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4399w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4405w4708w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4405w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4411w4716w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4411w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4417w4724w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4417w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4421w4732w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4421w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4225w4740w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4225w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4267w4524w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4267w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4230w4748w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4230w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4232w4756w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4232w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4234w4764w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4234w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4236w4772w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4236w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4273w4532w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4273w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4279w4540w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4279w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4285w4548w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4285w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4291w4556w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4291w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4297w4564w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4297w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4303w4572w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4303w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4309w4580w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4309w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5092w5333w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5092w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5151w5415w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5151w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5157w5423w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5157w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5163w5431w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5163w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5169w5439w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5169w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5175w5447w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5175w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5181w5455w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5181w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5187w5463w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5187w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5193w5471w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5193w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5199w5479w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5199w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5205w5487w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5205w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5097w5343w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5097w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5211w5495w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5211w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5217w5503w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5217w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5223w5511w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5223w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5229w5519w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5229w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5235w5527w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5235w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5241w5535w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5241w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5247w5543w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5247w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5251w5551w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5251w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5057w5559w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5057w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5062w5567w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5062w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5103w5351w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5103w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5064w5575w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5064w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5066w5583w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5066w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5068w5591w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5068w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5070w5599w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5070w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5109w5359w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5109w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5115w5367w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5115w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5121w5375w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5121w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5127w5383w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5127w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5133w5391w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5133w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5139w5399w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5139w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5145w5407w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range5145w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5923w6155w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5923w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5982w6237w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5982w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5988w6245w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5988w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5994w6253w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5994w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6000w6261w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6000w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6006w6269w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6006w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6012w6277w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6012w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6018w6285w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6018w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6024w6293w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6024w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6030w6301w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6030w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6036w6309w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6036w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5928w6165w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5928w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6042w6317w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6042w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6048w6325w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6048w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6054w6333w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6054w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6060w6341w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6060w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6066w6349w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6066w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6072w6357w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6072w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6076w6365w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range6076w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5884w6373w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5884w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5889w6381w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5889w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5891w6389w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5891w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5934w6173w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5934w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5893w6397w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5893w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5895w6405w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5895w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5897w6413w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5897w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5899w6421w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5899w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5940w6181w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5940w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5946w6189w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5946w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5952w6197w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5952w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5958w6205w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5958w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5964w6213w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5964w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5970w6221w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5970w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5976w6229w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5976w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6749w6972w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6749w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6808w7054w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6808w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6814w7062w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6814w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6820w7070w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6820w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6826w7078w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6826w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6832w7086w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6832w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6838w7094w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6838w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6844w7102w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6844w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6850w7110w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6850w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6856w7118w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6856w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6862w7126w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6862w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6754w6982w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6754w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6868w7134w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6868w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6874w7142w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6874w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6880w7150w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6880w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6886w7158w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6886w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6892w7166w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6892w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6896w7174w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6896w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6706w7182w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6706w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6711w7190w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6711w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6713w7198w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6713w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6715w7206w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6715w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6760w6990w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6760w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6717w7214w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6717w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6719w7222w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6719w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6721w7230w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6721w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6723w7238w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6723w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6766w6998w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6766w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6772w7006w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6772w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6778w7014w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6778w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6784w7022w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6784w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6790w7030w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6790w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6796w7038w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6796w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6802w7046w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6802w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7714w7782w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7714w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7743w7865w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7743w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7746w7873w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7746w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7749w7881w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7749w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7752w7889w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7752w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7755w7897w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7755w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7758w7905w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7758w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7761w7913w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7761w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7764w7921w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7764w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7767w7929w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7767w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7770w7937w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7770w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7716w7793w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7716w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7773w7945w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7773w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7776w7953w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7776w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7779w7961w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7779w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7544w7969w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7544w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7548w7977w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7548w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7550w7985w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7550w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7552w7993w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7552w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7554w8001w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7554w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7556w8009w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7556w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7558w8017w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7558w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7719w7801w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7719w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7560w8025w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7560w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7562w8033w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7562w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7564w8041w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7564w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7566w8049w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7566w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7722w7809w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7722w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7725w7817w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7725w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7728w7825w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7728w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7731w7833w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7731w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7734w7841w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7734w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7737w7849w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7737w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7740w7857w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7740w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8524w8589w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8524w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8553w8672w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8553w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8556w8680w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8556w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8559w8688w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8559w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8562w8696w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8562w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8565w8704w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8565w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8568w8712w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8568w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8571w8720w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8571w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8574w8728w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8574w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8577w8736w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8577w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8580w8744w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8580w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8526w8600w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8526w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8583w8752w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8583w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8586w8760w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8586w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8358w8768w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8358w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8362w8776w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8362w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8364w8784w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8364w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8366w8792w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8366w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8368w8800w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8368w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8370w8808w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8370w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8372w8816w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8372w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8374w8824w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8374w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8529w8608w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8529w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8376w8832w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8376w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8378w8840w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8378w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8380w8848w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8380w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8382w8856w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8382w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8532w8616w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8532w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8535w8624w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8535w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8538w8632w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8538w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8541w8640w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8541w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8544w8648w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8544w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8547w8656w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8547w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8550w8664w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8550w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9329w9391w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9329w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9358w9474w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9358w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9361w9482w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9361w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9364w9490w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9364w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9367w9498w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9367w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9370w9506w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9370w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9373w9514w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9373w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9376w9522w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9376w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9379w9530w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9379w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9382w9538w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9382w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9385w9546w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9385w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9331w9402w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9331w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9388w9554w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9388w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9167w9562w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9167w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9171w9570w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9171w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9173w9578w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9173w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9175w9586w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9175w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9177w9594w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9177w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9179w9602w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9179w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9181w9610w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9181w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9183w9618w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9183w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9185w9626w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9185w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9334w9410w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9334w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9187w9634w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9187w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9189w9642w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9189w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9191w9650w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9191w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9193w9658w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9193w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9337w9418w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9337w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9340w9426w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9340w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9343w9434w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9343w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9346w9442w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9346w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9349w9450w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9349w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9352w9458w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9352w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9355w9466w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9355w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10129w10188w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10129w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10158w10271w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10158w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10161w10279w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10161w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10164w10287w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10164w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10167w10295w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10167w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10170w10303w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10170w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10173w10311w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10173w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10176w10319w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10176w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10179w10327w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10179w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10182w10335w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10182w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10185w10343w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10185w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10131w10199w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10131w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9971w10351w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9971w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9975w10359w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9975w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9977w10367w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9977w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9979w10375w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9979w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9981w10383w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9981w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9983w10391w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9983w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9985w10399w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9985w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9987w10407w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9987w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9989w10415w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9989w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9991w10423w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9991w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10134w10207w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10134w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9993w10431w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9993w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9995w10439w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9995w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9997w10447w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9997w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9999w10455w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9999w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10137w10215w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10137w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10140w10223w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10140w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10143w10231w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10143w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10146w10239w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10146w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10149w10247w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10149w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10152w10255w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10152w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10155w10263w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10155w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1054w1146w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1054w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1083w1229w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1083w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1086w1237w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1086w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1089w1245w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1089w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1092w1253w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1092w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1095w1261w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1095w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1098w1269w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1098w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1101w1277w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1101w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1104w1285w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1104w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1107w1293w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1107w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1110w1301w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1110w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1056w1157w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1056w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1113w1309w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1113w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1116w1317w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1116w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1119w1325w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1119w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1122w1333w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1122w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1125w1341w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1125w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1128w1349w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1128w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1131w1357w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1131w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1134w1365w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1134w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1137w1373w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1137w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1140w1381w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1140w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1059w1165w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1059w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1143w1389w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1143w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range852w1397w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range852w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range856w1405w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range856w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range858w1413w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range858w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1062w1173w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1062w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1065w1181w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1065w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1068w1189w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1068w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1071w1197w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1071w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1074w1205w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1074w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1077w1213w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1077w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1080w1221w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1080w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1904w1993w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1904w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1933w2076w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1933w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1936w2084w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1936w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1939w2092w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1939w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1942w2100w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1942w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1945w2108w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1945w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1948w2116w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1948w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1951w2124w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1951w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1954w2132w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1954w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1957w2140w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1957w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1960w2148w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1960w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1906w2004w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1906w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1963w2156w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1963w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1966w2164w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1966w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1969w2172w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1969w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1972w2180w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1972w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1975w2188w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1975w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1978w2196w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1978w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1981w2204w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1981w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1984w2212w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1984w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1987w2220w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1987w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1990w2228w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1990w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1909w2012w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1909w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1706w2236w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1706w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1710w2244w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1710w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1712w2252w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1712w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1714w2260w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1714w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1912w2020w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1912w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1915w2028w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1915w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1918w2036w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1918w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1921w2044w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1921w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1924w2052w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1924w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1927w2060w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1927w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1930w2068w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1930w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2749w2835w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2749w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2778w2918w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2778w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2781w2926w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2781w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2784w2934w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2784w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2787w2942w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2787w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2790w2950w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2790w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2793w2958w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2793w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2796w2966w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2796w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2799w2974w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2799w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2802w2982w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2802w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2805w2990w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2805w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2751w2846w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2751w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2808w2998w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2808w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2811w3006w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2811w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2814w3014w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2814w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2817w3022w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2817w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2820w3030w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2820w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2823w3038w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2823w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2826w3046w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2826w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2829w3054w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2829w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2832w3062w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2832w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2555w3070w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2555w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2754w2854w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2754w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2559w3078w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2559w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2561w3086w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2561w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2563w3094w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2563w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2565w3102w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2565w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2757w2862w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2757w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2760w2870w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2760w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2763w2878w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2763w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2766w2886w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2766w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2769w2894w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2769w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2772w2902w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2772w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2775w2910w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2775w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3589w3672w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3589w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3618w3755w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3618w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3621w3763w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3621w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3624w3771w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3624w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3627w3779w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3627w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3630w3787w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3630w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3633w3795w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3633w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3636w3803w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3636w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3639w3811w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3639w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3642w3819w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3642w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3645w3827w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3645w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3591w3683w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3591w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3648w3835w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3648w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3651w3843w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3651w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3654w3851w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3654w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3657w3859w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3657w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3660w3867w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3660w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3663w3875w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3663w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3666w3883w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3666w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3669w3891w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3669w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3399w3899w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3399w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3403w3907w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3403w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3594w3691w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3594w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3405w3915w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3405w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3407w3923w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3407w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3409w3931w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3409w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3411w3939w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3411w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3597w3699w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3597w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3600w3707w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3600w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3603w3715w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3603w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3606w3723w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3606w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3609w3731w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3609w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3612w3739w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3612w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3615w3747w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3615w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4424w4504w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4424w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4453w4587w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4453w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4456w4595w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4456w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4459w4603w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4459w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4462w4611w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4462w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4465w4619w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4465w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4468w4627w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4468w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4471w4635w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4471w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4474w4643w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4474w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4477w4651w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4477w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4480w4659w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4480w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4426w4515w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4426w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4483w4667w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4483w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4486w4675w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4486w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4489w4683w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4489w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4492w4691w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4492w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4495w4699w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4495w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4498w4707w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4498w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4501w4715w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4501w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4238w4723w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4238w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4242w4731w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4242w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4244w4739w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4244w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4429w4523w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4429w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4246w4747w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4246w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4248w4755w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4248w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4250w4763w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4250w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4252w4771w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4252w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4432w4531w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4432w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4435w4539w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4435w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4438w4547w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4438w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4441w4555w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4441w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4444w4563w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4444w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4447w4571w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4447w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4450w4579w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4450w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5254w5331w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5254w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5283w5414w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5283w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5286w5422w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5286w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5289w5430w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5289w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5292w5438w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5292w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5295w5446w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5295w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5298w5454w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5298w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5301w5462w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5301w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5304w5470w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5304w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5307w5478w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5307w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5310w5486w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5310w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5256w5342w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5256w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5313w5494w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5313w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5316w5502w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5316w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5319w5510w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5319w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5322w5518w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5322w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5325w5526w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5325w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5328w5534w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5328w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5072w5542w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5072w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5076w5550w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5076w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5078w5558w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5078w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5080w5566w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5080w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5259w5350w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5259w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5082w5574w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5082w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5084w5582w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5084w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5086w5590w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5086w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5088w5598w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5088w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5262w5358w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5262w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5265w5366w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5265w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5268w5374w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5268w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5271w5382w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5271w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5274w5390w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5274w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5277w5398w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5277w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5280w5406w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5280w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6079w6153w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6079w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6108w6236w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6108w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6111w6244w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6111w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6114w6252w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6114w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6117w6260w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6117w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6120w6268w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6120w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6123w6276w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6123w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6126w6284w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6126w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6129w6292w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6129w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6132w6300w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6132w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6135w6308w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6135w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6081w6164w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6081w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6138w6316w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6138w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6141w6324w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6141w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6144w6332w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6144w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6147w6340w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6147w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6150w6348w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6150w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5901w6356w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5901w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5905w6364w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5905w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5907w6372w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5907w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5909w6380w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5909w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5911w6388w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5911w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6084w6172w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6084w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5913w6396w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5913w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5915w6404w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5915w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5917w6412w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5917w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5919w6420w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5919w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6087w6180w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6087w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6090w6188w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6090w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6093w6196w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6093w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6096w6204w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6096w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6099w6212w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6099w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6102w6220w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6102w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6105w6228w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6105w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6899w6970w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6899w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6928w7053w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6928w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6931w7061w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6931w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6934w7069w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6934w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6937w7077w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6937w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6940w7085w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6940w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6943w7093w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6943w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6946w7101w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6946w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6949w7109w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6949w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6952w7117w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6952w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6955w7125w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6955w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6901w6981w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6901w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6958w7133w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6958w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6961w7141w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6961w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6964w7149w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6964w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6967w7157w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6967w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6725w7165w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6725w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6729w7173w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6729w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6731w7181w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6731w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6733w7189w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6733w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6735w7197w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6735w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6737w7205w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6737w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6904w6989w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6904w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6739w7213w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6739w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6741w7221w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6741w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6743w7229w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6743w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6745w7237w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6745w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6907w6997w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6907w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6910w7005w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6910w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6913w7013w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6913w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6916w7021w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6916w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6919w7029w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6919w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6922w7037w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6922w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6925w7045w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6925w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7572w7789w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7572w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7631w7870w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7631w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7637w7878w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7637w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7643w7886w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7643w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7649w7894w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7649w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7655w7902w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7655w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7661w7910w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7661w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7667w7918w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7667w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7673w7926w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7673w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7679w7934w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7679w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7685w7942w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7685w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7577w7798w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7577w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7691w7950w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7691w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7697w7958w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7697w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7703w7966w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7703w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7709w7974w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7709w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7712w7982w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7712w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7526w7990w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7526w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7529w7998w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7529w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7531w8006w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7531w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7533w8014w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7533w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7535w8022w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7535w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7583w7806w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7583w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7537w8030w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7537w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7539w8038w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7539w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7541w8046w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7541w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7543w8054w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7543w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7589w7814w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7589w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7595w7822w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7595w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7601w7830w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7601w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7607w7838w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7607w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7613w7846w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7613w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7619w7854w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7619w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7625w7862w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7625w(0) AND wire_indexbitff_w_lg_w_q_range607w7783w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8388w8596w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8388w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8447w8677w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8447w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8453w8685w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8453w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8459w8693w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8459w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8465w8701w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8465w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8471w8709w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8471w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8477w8717w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8477w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8483w8725w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8483w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8489w8733w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8489w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8495w8741w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8495w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8501w8749w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8501w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8393w8605w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8393w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8507w8757w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8507w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8513w8765w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8513w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8519w8773w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8519w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8522w8781w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8522w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8338w8789w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8338w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8341w8797w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8341w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8343w8805w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8343w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8345w8813w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8345w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8347w8821w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8347w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8349w8829w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8349w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8399w8613w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8399w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8351w8837w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8351w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8353w8845w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8353w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8355w8853w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8355w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8357w8861w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8357w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8405w8621w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8405w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8411w8629w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8411w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8417w8637w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8417w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8423w8645w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8423w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8429w8653w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8429w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8435w8661w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8435w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8441w8669w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range8441w(0) AND wire_indexbitff_w_lg_w_q_range610w8590w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9199w9398w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9199w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9258w9479w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9258w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9264w9487w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9264w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9270w9495w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9270w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9276w9503w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9276w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9282w9511w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9282w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9288w9519w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9288w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9294w9527w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9294w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9300w9535w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9300w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9306w9543w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9306w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9312w9551w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9312w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9204w9407w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9204w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9318w9559w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9318w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9324w9567w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9324w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9327w9575w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9327w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9145w9583w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9145w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9148w9591w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9148w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9150w9599w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9150w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9152w9607w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9152w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9154w9615w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9154w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9156w9623w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9156w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9158w9631w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9158w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9210w9415w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9210w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9160w9639w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9160w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9162w9647w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9162w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9164w9655w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9164w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9166w9663w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9166w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9216w9423w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9216w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9222w9431w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9222w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9228w9439w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9228w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9234w9447w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9234w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9240w9455w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9240w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9246w9463w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9246w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9252w9471w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range9252w(0) AND wire_indexbitff_w_lg_w_q_range613w9392w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10005w10195w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10005w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10064w10276w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10064w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10070w10284w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10070w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10076w10292w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10076w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10082w10300w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10082w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10088w10308w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10088w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10094w10316w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10094w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10100w10324w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10100w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10106w10332w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10106w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10112w10340w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10112w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10118w10348w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10118w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10010w10204w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10010w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10124w10356w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10124w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10127w10364w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10127w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9947w10372w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9947w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9950w10380w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9950w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9952w10388w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9952w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9954w10396w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9954w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9956w10404w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9956w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9958w10412w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9958w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9960w10420w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9960w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9962w10428w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9962w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10016w10212w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10016w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9964w10436w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9964w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9966w10444w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9966w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9968w10452w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9968w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9970w10460w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9970w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10022w10220w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10022w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10028w10228w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10028w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10034w10236w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10034w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10040w10244w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10040w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10046w10252w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10046w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10052w10260w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10052w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10058w10268w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range10058w(0) AND wire_indexbitff_w_lg_w_q_range616w10189w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range864w1153w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range864w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range923w1234w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range923w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range929w1242w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range929w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range935w1250w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range935w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range941w1258w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range941w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range947w1266w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range947w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range953w1274w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range953w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range959w1282w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range959w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range965w1290w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range965w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range971w1298w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range971w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range977w1306w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range977w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range869w1162w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range869w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range983w1314w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range983w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range989w1322w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range989w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range995w1330w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range995w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1001w1338w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1001w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1007w1346w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1007w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1013w1354w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1013w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1019w1362w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1019w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1025w1370w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1025w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1031w1378w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1031w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1037w1386w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1037w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range875w1170w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range875w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1043w1394w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1043w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1049w1402w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1049w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1052w1410w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range1052w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range850w1418w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range850w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range881w1178w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range881w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range887w1186w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range887w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range893w1194w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range893w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range899w1202w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range899w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range905w1210w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range905w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range911w1218w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range911w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range917w1226w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range917w(0) AND wire_indexbitff_w_lg_w_q_range583w1147w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1720w2000w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1720w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1779w2081w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1779w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1785w2089w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1785w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1791w2097w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1791w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1797w2105w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1797w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1803w2113w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1803w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1809w2121w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1809w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1815w2129w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1815w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1821w2137w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1821w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1827w2145w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1827w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1833w2153w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1833w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1725w2009w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1725w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1839w2161w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1839w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1845w2169w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1845w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1851w2177w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1851w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1857w2185w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1857w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1863w2193w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1863w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1869w2201w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1869w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1875w2209w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1875w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1881w2217w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1881w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1887w2225w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1887w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1893w2233w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1893w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1731w2017w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1731w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1899w2241w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1899w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1902w2249w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1902w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1702w2257w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1702w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1705w2265w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1705w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1737w2025w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1737w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1743w2033w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1743w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1749w2041w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1749w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1755w2049w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1755w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1761w2057w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1761w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1767w2065w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1767w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1773w2073w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1773w(0) AND wire_indexbitff_w_lg_w_q_range586w1994w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2571w2842w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2571w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2630w2923w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2630w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2636w2931w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2636w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2642w2939w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2642w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2648w2947w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2648w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2654w2955w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2654w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2660w2963w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2660w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2666w2971w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2666w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2672w2979w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2672w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2678w2987w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2678w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2684w2995w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2684w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2576w2851w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2576w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2690w3003w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2690w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2696w3011w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2696w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2702w3019w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2702w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2708w3027w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2708w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2714w3035w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2714w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2720w3043w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2720w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2726w3051w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2726w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2732w3059w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2732w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2738w3067w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2738w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2744w3075w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2744w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2582w2859w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2582w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2747w3083w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2747w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2549w3091w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2549w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2552w3099w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2552w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2554w3107w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2554w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2588w2867w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2588w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2594w2875w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2594w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2600w2883w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2600w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2606w2891w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2606w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2612w2899w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2612w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2618w2907w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2618w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2624w2915w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2624w(0) AND wire_indexbitff_w_lg_w_q_range589w2836w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3417w3679w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3417w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3476w3760w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3476w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3482w3768w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3482w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3488w3776w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3488w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3494w3784w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3494w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3500w3792w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3500w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3506w3800w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3506w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3512w3808w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3512w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3518w3816w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3518w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3524w3824w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3524w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3530w3832w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3530w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3422w3688w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3422w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3536w3840w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3536w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3542w3848w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3542w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3548w3856w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3548w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3554w3864w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3554w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3560w3872w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3560w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3566w3880w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3566w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3572w3888w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3572w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3578w3896w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3578w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3584w3904w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3584w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3587w3912w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3587w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3428w3696w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3428w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3391w3920w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3391w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3394w3928w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3394w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3396w3936w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3396w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3398w3944w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3398w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3434w3704w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3434w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3440w3712w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3440w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3446w3720w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3446w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3452w3728w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3452w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3458w3736w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3458w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3464w3744w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3464w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3470w3752w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3470w(0) AND wire_indexbitff_w_lg_w_q_range592w3673w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4258w4511w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4258w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4317w4592w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4317w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4323w4600w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4323w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4329w4608w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4329w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4335w4616w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4335w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4341w4624w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4341w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4347w4632w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4347w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4353w4640w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4353w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4359w4648w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4359w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4365w4656w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4365w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4371w4664w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4371w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4263w4520w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4263w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4377w4672w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4377w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4383w4680w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4383w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4389w4688w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4389w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4395w4696w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4395w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4401w4704w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4401w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4407w4712w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4407w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4413w4720w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4413w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4419w4728w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4419w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4422w4736w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4422w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4228w4744w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4228w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4269w4528w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4269w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4231w4752w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4231w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4233w4760w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4233w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4235w4768w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4235w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4237w4776w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4237w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4275w4536w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4275w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4281w4544w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4281w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4287w4552w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4287w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4293w4560w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4293w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4299w4568w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4299w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4305w4576w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4305w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4311w4584w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4311w(0) AND wire_indexbitff_w_lg_w_q_range595w4505w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5094w5338w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5094w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5153w5419w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5153w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5159w5427w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5159w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5165w5435w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5165w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5171w5443w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5171w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5177w5451w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5177w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5183w5459w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5183w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5189w5467w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5189w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5195w5475w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5195w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5201w5483w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5201w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5207w5491w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5207w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5099w5347w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5099w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5213w5499w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5213w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5219w5507w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5219w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5225w5515w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5225w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5231w5523w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5231w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5237w5531w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5237w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5243w5539w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5243w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5249w5547w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5249w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5252w5555w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5252w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5060w5563w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5060w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5063w5571w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5063w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5105w5355w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5105w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5065w5579w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5065w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5067w5587w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5067w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5069w5595w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5069w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5071w5603w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5071w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5111w5363w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5111w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5117w5371w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5117w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5123w5379w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5123w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5129w5387w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5129w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5135w5395w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5135w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5141w5403w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5141w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5147w5411w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range5147w(0) AND wire_indexbitff_w_lg_w_q_range598w5332w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5925w6160w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5925w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5984w6241w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5984w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5990w6249w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5990w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5996w6257w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5996w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6002w6265w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6002w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6008w6273w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6008w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6014w6281w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6014w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6020w6289w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6020w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6026w6297w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6026w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6032w6305w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6032w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6038w6313w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6038w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5930w6169w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5930w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6044w6321w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6044w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6050w6329w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6050w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6056w6337w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6056w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6062w6345w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6062w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6068w6353w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6068w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6074w6361w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6074w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6077w6369w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range6077w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5887w6377w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5887w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5890w6385w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5890w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5892w6393w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5892w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5936w6177w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5936w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5894w6401w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5894w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5896w6409w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5896w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5898w6417w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5898w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5900w6425w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5900w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5942w6185w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5942w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5948w6193w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5948w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5954w6201w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5954w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5960w6209w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5960w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5966w6217w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5966w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5972w6225w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5972w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5978w6233w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5978w(0) AND wire_indexbitff_w_lg_w_q_range601w6154w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6751w6977w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6751w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6810w7058w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6810w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6816w7066w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6816w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6822w7074w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6822w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6828w7082w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6828w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6834w7090w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6834w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6840w7098w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6840w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6846w7106w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6846w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6852w7114w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6852w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6858w7122w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6858w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6864w7130w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6864w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6756w6986w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6756w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6870w7138w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6870w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6876w7146w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6876w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6882w7154w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6882w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6888w7162w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6888w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6894w7170w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6894w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6897w7178w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6897w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6709w7186w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6709w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6712w7194w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6712w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6714w7202w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6714w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6716w7210w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6716w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6762w6994w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6762w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6718w7218w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6718w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6720w7226w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6720w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6722w7234w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6722w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6724w7242w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6724w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6768w7002w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6768w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6774w7010w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6774w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6780w7018w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6780w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6786w7026w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6786w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6792w7034w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6792w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6798w7042w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6798w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6804w7050w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6804w(0) AND wire_indexbitff_w_lg_w_q_range604w6971w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7715w7788w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7715w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7744w7869w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7744w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7747w7877w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7747w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7750w7885w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7750w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7753w7893w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7753w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7756w7901w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7756w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7759w7909w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7759w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7762w7917w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7762w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7765w7925w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7765w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7768w7933w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7768w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7771w7941w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7771w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7717w7797w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7717w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7774w7949w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7774w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7777w7957w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7777w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7780w7965w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7780w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7546w7973w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7546w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7549w7981w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7549w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7551w7989w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7551w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7553w7997w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7553w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7555w8005w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7555w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7557w8013w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7557w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7559w8021w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7559w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7720w7805w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7720w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7561w8029w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7561w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7563w8037w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7563w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7565w8045w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7565w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7567w8053w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7567w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7723w7813w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7723w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7726w7821w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7726w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7729w7829w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7729w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7732w7837w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7732w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7735w7845w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7735w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7738w7853w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7738w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7741w7861w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7741w(0) AND wire_indexbitff_w_q_range607w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8525w8595w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8525w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8554w8676w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8554w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8557w8684w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8557w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8560w8692w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8560w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8563w8700w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8563w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8566w8708w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8566w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8569w8716w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8569w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8572w8724w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8572w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8575w8732w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8575w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8578w8740w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8578w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8581w8748w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8581w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8527w8604w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8527w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8584w8756w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8584w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8587w8764w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8587w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8360w8772w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8360w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8363w8780w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8363w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8365w8788w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8365w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8367w8796w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8367w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8369w8804w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8369w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8371w8812w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8371w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8373w8820w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8373w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8375w8828w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8375w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8530w8612w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8530w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8377w8836w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8377w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8379w8844w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8379w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8381w8852w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8381w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8383w8860w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8383w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8533w8620w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8533w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8536w8628w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8536w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8539w8636w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8539w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8542w8644w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8542w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8545w8652w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8545w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8548w8660w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8548w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8551w8668w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8551w(0) AND wire_indexbitff_w_q_range610w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9330w9397w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9330w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9359w9478w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9359w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9362w9486w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9362w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9365w9494w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9365w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9368w9502w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9368w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9371w9510w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9371w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9374w9518w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9374w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9377w9526w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9377w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9380w9534w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9380w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9383w9542w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9383w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9386w9550w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9386w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9332w9406w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9332w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9389w9558w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9389w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9169w9566w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9169w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9172w9574w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9172w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9174w9582w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9174w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9176w9590w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9176w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9178w9598w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9178w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9180w9606w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9180w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9182w9614w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9182w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9184w9622w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9184w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9186w9630w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9186w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9335w9414w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9335w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9188w9638w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9188w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9190w9646w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9190w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9192w9654w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9192w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9194w9662w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9194w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9338w9422w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9338w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9341w9430w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9341w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9344w9438w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9344w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9347w9446w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9347w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9350w9454w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9350w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9353w9462w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9353w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9356w9470w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9356w(0) AND wire_indexbitff_w_q_range613w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10130w10194w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10130w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10159w10275w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10159w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10162w10283w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10162w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10165w10291w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10165w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10168w10299w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10168w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10171w10307w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10171w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10174w10315w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10174w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10177w10323w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10177w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10180w10331w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10180w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10183w10339w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10183w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10186w10347w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10186w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10132w10203w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10132w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9973w10355w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9973w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9976w10363w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9976w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9978w10371w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9978w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9980w10379w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9980w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9982w10387w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9982w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9984w10395w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9984w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9986w10403w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9986w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9988w10411w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9988w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9990w10419w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9990w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9992w10427w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9992w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10135w10211w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10135w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9994w10435w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9994w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9996w10443w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9996w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9998w10451w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9998w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10000w10459w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10000w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10138w10219w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10138w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10141w10227w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10141w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10144w10235w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10144w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10147w10243w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10147w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10150w10251w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10150w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10153w10259w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10153w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10156w10267w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10156w(0) AND wire_indexbitff_w_q_range616w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1055w1152w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1055w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1084w1233w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1084w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1087w1241w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1087w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1090w1249w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1090w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1093w1257w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1093w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1096w1265w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1096w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1099w1273w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1099w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1102w1281w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1102w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1105w1289w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1105w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1108w1297w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1108w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1111w1305w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1111w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1057w1161w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1057w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1114w1313w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1114w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1117w1321w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1117w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1120w1329w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1120w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1123w1337w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1123w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1126w1345w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1126w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1129w1353w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1129w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1132w1361w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1132w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1135w1369w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1135w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1138w1377w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1138w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1141w1385w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1141w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1060w1169w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1060w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1144w1393w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1144w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range854w1401w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range854w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range857w1409w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range857w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range859w1417w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range859w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1063w1177w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1063w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1066w1185w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1066w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1069w1193w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1069w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1072w1201w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1072w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1075w1209w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1075w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1078w1217w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1078w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1081w1225w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1081w(0) AND wire_indexbitff_w_q_range583w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1905w1999w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1905w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1934w2080w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1934w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1937w2088w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1937w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1940w2096w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1940w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1943w2104w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1943w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1946w2112w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1946w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1949w2120w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1949w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1952w2128w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1952w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1955w2136w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1955w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1958w2144w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1958w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1961w2152w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1961w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1907w2008w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1907w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1964w2160w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1964w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1967w2168w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1967w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1970w2176w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1970w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1973w2184w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1973w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1976w2192w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1976w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1979w2200w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1979w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1982w2208w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1982w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1985w2216w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1985w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1988w2224w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1988w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1991w2232w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1991w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1910w2016w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1910w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1708w2240w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1708w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1711w2248w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1711w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1713w2256w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1713w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1715w2264w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1715w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1913w2024w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1913w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1916w2032w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1916w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1919w2040w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1919w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1922w2048w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1922w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1925w2056w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1925w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1928w2064w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1928w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1931w2072w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1931w(0) AND wire_indexbitff_w_q_range586w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2750w2841w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2750w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2779w2922w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2779w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2782w2930w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2782w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2785w2938w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2785w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2788w2946w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2788w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2791w2954w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2791w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2794w2962w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2794w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2797w2970w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2797w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2800w2978w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2800w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2803w2986w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2803w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2806w2994w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2806w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2752w2850w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2752w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2809w3002w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2809w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2812w3010w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2812w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2815w3018w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2815w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2818w3026w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2818w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2821w3034w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2821w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2824w3042w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2824w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2827w3050w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2827w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2830w3058w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2830w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2833w3066w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2833w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2557w3074w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2557w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2755w2858w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2755w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2560w3082w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2560w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2562w3090w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2562w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2564w3098w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2564w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2566w3106w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2566w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2758w2866w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2758w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2761w2874w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2761w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2764w2882w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2764w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2767w2890w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2767w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2770w2898w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2770w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2773w2906w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2773w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2776w2914w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2776w(0) AND wire_indexbitff_w_q_range589w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3590w3678w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3590w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3619w3759w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3619w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3622w3767w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3622w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3625w3775w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3625w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3628w3783w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3628w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3631w3791w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3631w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3634w3799w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3634w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3637w3807w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3637w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3640w3815w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3640w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3643w3823w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3643w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3646w3831w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3646w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3592w3687w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3592w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3649w3839w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3649w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3652w3847w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3652w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3655w3855w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3655w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3658w3863w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3658w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3661w3871w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3661w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3664w3879w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3664w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3667w3887w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3667w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3670w3895w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3670w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3401w3903w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3401w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3404w3911w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3404w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3595w3695w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3595w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3406w3919w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3406w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3408w3927w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3408w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3410w3935w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3410w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3412w3943w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3412w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3598w3703w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3598w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3601w3711w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3601w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3604w3719w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3604w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3607w3727w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3607w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3610w3735w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3610w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3613w3743w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3613w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3616w3751w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3616w(0) AND wire_indexbitff_w_q_range592w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4425w4510w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4425w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4454w4591w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4454w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4457w4599w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4457w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4460w4607w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4460w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4463w4615w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4463w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4466w4623w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4466w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4469w4631w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4469w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4472w4639w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4472w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4475w4647w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4475w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4478w4655w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4478w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4481w4663w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4481w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4427w4519w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4427w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4484w4671w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4484w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4487w4679w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4487w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4490w4687w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4490w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4493w4695w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4493w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4496w4703w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4496w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4499w4711w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4499w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4502w4719w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4502w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4240w4727w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4240w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4243w4735w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4243w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4245w4743w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4245w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4430w4527w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4430w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4247w4751w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4247w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4249w4759w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4249w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4251w4767w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4251w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4253w4775w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4253w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4433w4535w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4433w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4436w4543w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4436w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4439w4551w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4439w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4442w4559w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4442w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4445w4567w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4445w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4448w4575w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4448w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4451w4583w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4451w(0) AND wire_indexbitff_w_q_range595w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5255w5337w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5255w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5284w5418w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5284w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5287w5426w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5287w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5290w5434w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5290w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5293w5442w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5293w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5296w5450w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5296w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5299w5458w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5299w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5302w5466w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5302w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5305w5474w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5305w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5308w5482w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5308w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5311w5490w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5311w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5257w5346w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5257w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5314w5498w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5314w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5317w5506w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5317w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5320w5514w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5320w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5323w5522w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5323w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5326w5530w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5326w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5329w5538w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5329w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5074w5546w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5074w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5077w5554w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5077w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5079w5562w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5079w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5081w5570w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5081w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5260w5354w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5260w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5083w5578w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5083w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5085w5586w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5085w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5087w5594w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5087w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5089w5602w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5089w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5263w5362w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5263w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5266w5370w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5266w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5269w5378w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5269w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5272w5386w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5272w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5275w5394w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5275w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5278w5402w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5278w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5281w5410w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5281w(0) AND wire_indexbitff_w_q_range598w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6080w6159w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6080w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6109w6240w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6109w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6112w6248w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6112w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6115w6256w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6115w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6118w6264w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6118w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6121w6272w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6121w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6124w6280w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6124w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6127w6288w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6127w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6130w6296w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6130w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6133w6304w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6133w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6136w6312w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6136w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6082w6168w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6082w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6139w6320w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6139w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6142w6328w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6142w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6145w6336w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6145w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6148w6344w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6148w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6151w6352w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6151w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5903w6360w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5903w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5906w6368w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5906w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5908w6376w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5908w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5910w6384w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5910w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5912w6392w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5912w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6085w6176w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6085w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5914w6400w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5914w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5916w6408w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5916w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5918w6416w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5918w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5920w6424w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5920w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6088w6184w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6088w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6091w6192w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6091w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6094w6200w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6094w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6097w6208w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6097w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6100w6216w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6100w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6103w6224w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6103w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6106w6232w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6106w(0) AND wire_indexbitff_w_q_range601w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6900w6976w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6900w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6929w7057w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6929w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6932w7065w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6932w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6935w7073w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6935w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6938w7081w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6938w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6941w7089w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6941w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6944w7097w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6944w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6947w7105w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6947w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6950w7113w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6950w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6953w7121w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6953w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6956w7129w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6956w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6902w6985w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6902w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6959w7137w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6959w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6962w7145w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6962w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6965w7153w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6965w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6968w7161w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6968w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6727w7169w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6727w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6730w7177w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6730w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6732w7185w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6732w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6734w7193w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6734w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6736w7201w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6736w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6738w7209w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6738w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6905w6993w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6905w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6740w7217w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6740w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6742w7225w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6742w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6744w7233w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6744w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6746w7241w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6746w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6908w7001w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6908w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6911w7009w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6911w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6914w7017w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6914w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6917w7025w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6917w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6920w7033w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6920w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6923w7041w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6923w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6926w7049w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6926w(0) AND wire_indexbitff_w_q_range604w(0);
	wire_ccc_cordic_m_w_lg_indexbit412w(0) <= NOT indexbit;
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8871w8872w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8871w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8952w8953w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8952w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8960w8961w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8960w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8968w8969w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8968w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8976w8977w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8984w8985w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8984w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8992w8993w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8992w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9000w9001w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9000w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9008w9009w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9008w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9016w9017w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9016w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9024w9025w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9024w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8880w8881w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8880w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9032w9033w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9032w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9040w9041w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9040w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9048w9049w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9048w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9056w9057w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9056w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9064w9065w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9064w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9072w9073w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9072w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9080w9081w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9080w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9088w9089w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9088w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9096w9097w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9096w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9104w9105w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9104w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8888w8889w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8888w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9112w9113w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9112w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9120w9121w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9120w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9128w9129w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9128w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9136w9137w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range9136w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8896w8897w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8896w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8904w8905w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8904w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8912w8913w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8912w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8920w8921w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8920w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8928w8929w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8928w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8936w8937w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8936w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8944w8945w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8944w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9673w9674w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9673w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9754w9755w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9754w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9762w9763w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9762w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9770w9771w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9770w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9778w9779w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9778w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9786w9787w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9786w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9794w9795w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9794w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9802w9803w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9802w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9810w9811w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9810w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9818w9819w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9818w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9826w9827w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9826w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9682w9683w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9682w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9834w9835w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9834w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9842w9843w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9842w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9850w9851w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9850w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9858w9859w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9858w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9866w9867w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9866w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9874w9875w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9874w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9882w9883w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9882w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9890w9891w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9890w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9898w9899w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9898w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9906w9907w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9906w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9690w9691w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9690w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9914w9915w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9914w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9922w9923w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9922w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9930w9931w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9930w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9938w9939w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9938w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9698w9699w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9698w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9706w9707w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9706w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9714w9715w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9714w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9722w9723w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9730w9731w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9730w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9738w9739w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9738w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9746w9747w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9746w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10470w10471w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10470w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10551w10552w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10551w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10559w10560w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10559w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10567w10568w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10567w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10575w10576w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10575w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10583w10584w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10583w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10591w10592w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10591w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10599w10600w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10599w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10607w10608w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10607w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10615w10616w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10615w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10623w10624w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10623w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10479w10480w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10479w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10631w10632w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10631w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10639w10640w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10639w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10647w10648w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10647w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10655w10656w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10655w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10663w10664w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10663w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10671w10672w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10671w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10679w10680w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10679w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10687w10688w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10687w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10695w10696w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10695w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10703w10704w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10703w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10487w10488w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10487w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10711w10712w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10711w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10719w10720w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10719w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10727w10728w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10727w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10735w10736w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10735w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10495w10496w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10495w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10503w10504w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10503w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10511w10512w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10511w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10519w10520w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10519w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10527w10528w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10527w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10535w10536w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10535w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10543w10544w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range10543w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1428w1429w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1428w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1509w1510w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1509w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1517w1518w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1517w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1525w1526w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1525w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1533w1534w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1533w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1541w1542w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1541w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1549w1550w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1549w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1557w1558w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1557w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1565w1566w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1565w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1573w1574w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1573w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1581w1582w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1581w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1437w1438w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1437w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1589w1590w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1589w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1597w1598w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1597w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1605w1606w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1605w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1613w1614w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1613w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1621w1622w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1621w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1629w1630w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1629w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1637w1638w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1637w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1645w1646w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1645w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1653w1654w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1653w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1661w1662w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1661w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1445w1446w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1445w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1669w1670w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1669w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1677w1678w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1677w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1685w1686w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1685w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1693w1694w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1693w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1453w1454w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1453w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1461w1462w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1461w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1469w1470w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1469w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1477w1478w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1477w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1485w1486w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1485w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1493w1494w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1493w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1501w1502w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1501w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2275w2276w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2275w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2356w2357w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2356w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2364w2365w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2364w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2372w2373w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2372w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2380w2381w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2380w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2388w2389w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2388w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2396w2397w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2396w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2404w2405w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2404w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2412w2413w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2412w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2420w2421w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2420w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2428w2429w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2428w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2284w2285w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2284w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2436w2437w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2436w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2444w2445w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2444w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2452w2453w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2452w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2460w2461w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2460w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2468w2469w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2468w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2476w2477w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2476w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2484w2485w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2484w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2492w2493w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2492w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2500w2501w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2500w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2508w2509w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2508w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2292w2293w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2292w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2516w2517w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2516w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2524w2525w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2524w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2532w2533w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2532w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2540w2541w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2540w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2300w2301w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2300w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2308w2309w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2308w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2316w2317w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2316w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2324w2325w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2324w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2332w2333w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2332w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2340w2341w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2340w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2348w2349w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2348w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3117w3118w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3117w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3198w3199w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3198w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3206w3207w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3206w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3214w3215w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3214w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3222w3223w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3222w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3230w3231w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3230w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3238w3239w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3238w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3246w3247w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3246w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3254w3255w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3254w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3262w3263w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3262w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3270w3271w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3270w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3126w3127w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3126w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3278w3279w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3278w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3286w3287w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3286w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3294w3295w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3294w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3302w3303w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3302w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3310w3311w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3310w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3318w3319w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3318w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3326w3327w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3326w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3334w3335w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3334w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3342w3343w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3342w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3350w3351w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3350w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3134w3135w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3134w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3358w3359w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3358w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3366w3367w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3366w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3374w3375w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3374w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3382w3383w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3382w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3142w3143w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3142w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3150w3151w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3150w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3158w3159w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3158w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3166w3167w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3166w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3174w3175w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3174w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3182w3183w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3182w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3190w3191w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3190w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3954w3955w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3954w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4035w4036w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4035w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4043w4044w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4043w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4051w4052w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4051w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4059w4060w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4059w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4067w4068w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4067w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4075w4076w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4075w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4083w4084w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4083w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4091w4092w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4091w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4099w4100w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4099w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4107w4108w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4107w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3963w3964w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3963w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4115w4116w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4115w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4123w4124w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4123w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4131w4132w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4131w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4139w4140w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4139w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4147w4148w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4147w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4155w4156w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4155w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4163w4164w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4163w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4171w4172w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4171w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4179w4180w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4179w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4187w4188w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4187w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3971w3972w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3971w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4195w4196w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4195w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4203w4204w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4203w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4211w4212w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4211w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4219w4220w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4219w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3979w3980w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3979w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3987w3988w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3987w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3995w3996w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3995w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4003w4004w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4003w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4011w4012w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4011w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4019w4020w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4019w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4027w4028w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range4027w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4786w4787w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4786w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4867w4868w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4867w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4875w4876w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4875w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4883w4884w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4883w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4891w4892w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4891w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4899w4900w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4899w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4907w4908w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4907w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4915w4916w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4915w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4923w4924w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4923w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4931w4932w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4931w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4939w4940w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4939w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4795w4796w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4795w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4947w4948w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4947w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4955w4956w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4955w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4963w4964w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4963w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4971w4972w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4971w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4979w4980w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4979w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4987w4988w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4987w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4995w4996w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4995w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5003w5004w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5003w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5011w5012w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5011w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5019w5020w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5019w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4803w4804w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4803w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5027w5028w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5027w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5035w5036w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5035w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5043w5044w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5043w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5051w5052w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range5051w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4811w4812w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4811w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4819w4820w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4819w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4827w4828w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4827w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4835w4836w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4835w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4843w4844w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4843w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4851w4852w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4851w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4859w4860w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4859w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5613w5614w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5613w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5694w5695w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5694w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5702w5703w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5702w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5710w5711w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5710w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5718w5719w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5718w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5726w5727w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5726w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5734w5735w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5734w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5742w5743w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5742w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5750w5751w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5750w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5758w5759w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5758w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5766w5767w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5766w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5622w5623w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5622w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5774w5775w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5774w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5782w5783w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5782w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5790w5791w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5790w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5798w5799w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5798w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5806w5807w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5806w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5814w5815w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5814w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5822w5823w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5822w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5830w5831w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5830w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5838w5839w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5838w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5846w5847w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5846w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5630w5631w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5630w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5854w5855w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5854w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5862w5863w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5862w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5870w5871w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5870w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5878w5879w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5878w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5638w5639w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5638w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5646w5647w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5646w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5654w5655w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5654w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5662w5663w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5662w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5670w5671w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5670w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5678w5679w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5678w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5686w5687w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5686w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6435w6436w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6435w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6516w6517w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6516w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6524w6525w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6524w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6532w6533w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6532w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6540w6541w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6540w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6548w6549w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6548w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6556w6557w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6556w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6564w6565w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6564w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6572w6573w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6572w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6580w6581w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6580w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6588w6589w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6588w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6444w6445w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6444w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6596w6597w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6596w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6604w6605w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6604w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6612w6613w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6612w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6620w6621w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6620w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6628w6629w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6628w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6636w6637w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6636w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6644w6645w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6644w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6652w6653w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6652w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6660w6661w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6660w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6668w6669w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6668w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6452w6453w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6452w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6676w6677w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6676w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6684w6685w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6684w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6692w6693w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6692w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6700w6701w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6700w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6460w6461w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6460w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6468w6469w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6468w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6476w6477w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6476w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6484w6485w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6484w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6492w6493w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6492w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6500w6501w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6500w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6508w6509w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6508w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7252w7253w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7252w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7333w7334w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7333w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7341w7342w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7341w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7349w7350w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7349w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7357w7358w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7357w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7365w7366w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7365w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7373w7374w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7373w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7381w7382w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7381w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7389w7390w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7389w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7397w7398w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7397w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7405w7406w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7405w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7261w7262w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7261w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7413w7414w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7413w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7421w7422w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7421w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7429w7430w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7429w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7437w7438w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7437w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7445w7446w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7445w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7453w7454w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7453w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7461w7462w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7461w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7469w7470w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7477w7478w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7477w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7485w7486w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7485w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7269w7270w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7269w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7493w7494w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7493w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7501w7502w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7501w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7509w7510w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7509w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7517w7518w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7517w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7277w7278w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7277w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7285w7286w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7285w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7293w7294w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7293w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7301w7302w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7301w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7309w7310w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7309w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7317w7318w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7317w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7325w7326w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range7325w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8064w8065w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8064w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8145w8146w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8145w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8153w8154w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8153w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8161w8162w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8161w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8169w8170w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8169w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8177w8178w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8177w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8185w8186w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8185w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8193w8194w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8193w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8201w8202w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8201w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8209w8210w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8209w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8217w8218w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8217w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8073w8074w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8073w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8225w8226w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8233w8234w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8233w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8241w8242w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8241w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8249w8250w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8249w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8257w8258w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8257w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8265w8266w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8265w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8273w8274w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8273w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8281w8282w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8281w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8289w8290w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8289w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8297w8298w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8297w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8081w8082w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8081w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8305w8306w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8305w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8313w8314w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8313w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8321w8322w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8321w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8329w8330w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8329w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8089w8090w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8089w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8097w8098w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8097w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8105w8106w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8105w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8113w8114w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8113w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8121w8122w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8121w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8129w8130w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8129w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8137w8138w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range8137w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10753w10754w10755w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10753w10754w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10750w10751w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10794w10806w10807w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10794w10806w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10804w10805w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10799w10811w10812w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10799w10811w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10809w10810w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10804w10816w10817w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10804w10816w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10814w10815w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10809w10821w10822w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10809w10821w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10819w10820w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10814w10826w10827w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10814w10826w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10824w10825w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10819w10831w10832w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10819w10831w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10829w10830w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10824w10836w10837w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10824w10836w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10834w10835w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10829w10841w10842w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10829w10841w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10839w10840w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10834w10846w10847w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10834w10846w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10844w10845w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10839w10851w10852w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10839w10851w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10849w10850w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10760w10761w10762w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10760w10761w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10758w10759w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10844w10856w10857w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10844w10856w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10854w10855w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10849w10861w10862w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10849w10861w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10859w10860w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10854w10866w10867w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10854w10866w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10864w10865w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10859w10871w10872w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10859w10871w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10869w10870w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10864w10876w10877w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10864w10876w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10874w10875w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10869w10881w10882w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10869w10881w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10879w10880w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10874w10886w10887w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10874w10886w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10884w10885w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10879w10891w10892w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10879w10891w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10889w10890w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10884w10896w10897w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10884w10896w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10894w10895w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10889w10901w10902w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10889w10901w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10899w10900w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10750w10766w10767w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10750w10766w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10764w10765w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10894w10906w10907w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10894w10906w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10904w10905w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10899w10911w10912w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10899w10911w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10910w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10904w10914w10915w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10904w10914w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10910w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10909w10917w10918w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10917w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10909w10910w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10758w10771w10772w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10758w10771w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10769w10770w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10764w10776w10777w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10764w10776w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10774w10775w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10769w10781w10782w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10769w10781w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10779w10780w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10774w10786w10787w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10774w10786w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10784w10785w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10779w10791w10792w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10779w10791w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10789w10790w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10784w10796w10797w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10784w10796w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10794w10795w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10789w10801w10802w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10789w10801w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10799w10800w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range458w461w462w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range458w461w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range448w460w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range463w466w467w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range463w466w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range453w465w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range468w471w472w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range468w471w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range458w470w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range473w476w477w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range473w476w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range463w475w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range478w481w482w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range478w481w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range468w480w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range483w486w487w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range483w486w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range473w485w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range488w491w492w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range488w491w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range478w490w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range493w496w497w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range493w496w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range483w495w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range498w501w502w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range498w501w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range488w500w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range503w506w507w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range503w506w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range493w505w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range508w511w512w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range508w511w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range498w510w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range513w516w517w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range513w516w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range503w515w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range518w521w522w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range518w521w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range508w520w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range523w526w527w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range523w526w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range513w525w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range528w531w532w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range528w531w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range518w530w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range533w536w537w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range533w536w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range523w535w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range538w541w542w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range538w541w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range528w540w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range543w546w547w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range543w546w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range533w545w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range548w551w552w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range548w551w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range538w550w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range553w556w557w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range553w556w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range543w555w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range418w421w422w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range418w421w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range410w420w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range558w561w562w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range558w561w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range548w560w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range563w566w567w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range563w566w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range553w565w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range568w571w572w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range568w571w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range558w570w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range573w576w577w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range573w576w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range563w575w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range423w426w427w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range423w426w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range415w425w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range428w431w432w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range428w431w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range418w430w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range433w436w437w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range433w436w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range423w435w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range438w441w442w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range438w441w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range428w440w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range443w446w447w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range443w446w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range433w445w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range448w451w452w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range448w451w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range438w450w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range453w456w457w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range453w456w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range443w455w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7570w7784w7785w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7570w7784w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7714w7782w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7629w7866w7867w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7629w7866w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7743w7865w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7635w7874w7875w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7635w7874w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7746w7873w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7641w7882w7883w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7641w7882w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7749w7881w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7647w7890w7891w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7647w7890w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7752w7889w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7653w7898w7899w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7653w7898w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7755w7897w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7659w7906w7907w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7659w7906w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7758w7905w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7665w7914w7915w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7665w7914w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7761w7913w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7671w7922w7923w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7671w7922w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7764w7921w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7677w7930w7931w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7677w7930w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7767w7929w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7683w7938w7939w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7683w7938w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7770w7937w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7575w7794w7795w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7575w7794w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7716w7793w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7689w7946w7947w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7689w7946w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7773w7945w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7695w7954w7955w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7695w7954w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7776w7953w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7701w7962w7963w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7701w7962w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7779w7961w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7707w7970w7971w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7707w7970w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7544w7969w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7711w7978w7979w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7711w7978w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7548w7977w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7523w7986w7987w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7523w7986w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7550w7985w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7528w7994w7995w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7528w7994w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7552w7993w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7530w8002w8003w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7530w8002w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7554w8001w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7532w8010w8011w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7532w8010w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7556w8009w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7534w8018w8019w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7534w8018w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7558w8017w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7581w7802w7803w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7581w7802w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7719w7801w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7536w8026w8027w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7536w8026w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7560w8025w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7538w8034w8035w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7538w8034w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7562w8033w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7540w8042w8043w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7540w8042w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7564w8041w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7542w8050w8051w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7542w8050w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7566w8049w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7587w7810w7811w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7587w7810w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7722w7809w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7593w7818w7819w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7593w7818w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7725w7817w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7599w7826w7827w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7599w7826w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7728w7825w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7605w7834w7835w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7605w7834w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7731w7833w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7611w7842w7843w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7611w7842w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7734w7841w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7617w7850w7851w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7617w7850w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7737w7849w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7623w7858w7859w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7623w7858w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7740w7857w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8386w8591w8592w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8386w8591w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8524w8589w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8445w8673w8674w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8445w8673w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8553w8672w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8451w8681w8682w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8451w8681w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8556w8680w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8457w8689w8690w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8457w8689w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8559w8688w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8463w8697w8698w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8463w8697w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8562w8696w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8469w8705w8706w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8469w8705w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8565w8704w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8475w8713w8714w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8475w8713w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8568w8712w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8481w8721w8722w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8481w8721w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8571w8720w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8487w8729w8730w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8487w8729w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8574w8728w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8493w8737w8738w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8493w8737w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8577w8736w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8499w8745w8746w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8499w8745w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8580w8744w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8391w8601w8602w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8391w8601w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8526w8600w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8505w8753w8754w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8505w8753w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8583w8752w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8511w8761w8762w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8511w8761w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8586w8760w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8517w8769w8770w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8517w8769w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8358w8768w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8521w8777w8778w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8521w8777w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8362w8776w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8335w8785w8786w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8335w8785w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8364w8784w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8340w8793w8794w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8340w8793w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8366w8792w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8342w8801w8802w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8342w8801w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8368w8800w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8344w8809w8810w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8344w8809w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8370w8808w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8346w8817w8818w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8346w8817w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8372w8816w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8348w8825w8826w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8348w8825w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8374w8824w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8397w8609w8610w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8397w8609w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8529w8608w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8350w8833w8834w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8350w8833w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8376w8832w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8352w8841w8842w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8352w8841w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8378w8840w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8354w8849w8850w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8354w8849w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8380w8848w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8356w8857w8858w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8356w8857w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8382w8856w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8403w8617w8618w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8403w8617w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8532w8616w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8409w8625w8626w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8409w8625w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8535w8624w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8415w8633w8634w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8415w8633w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8538w8632w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8421w8641w8642w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8421w8641w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8541w8640w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8427w8649w8650w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8427w8649w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8544w8648w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8433w8657w8658w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8433w8657w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8547w8656w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8439w8665w8666w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range8439w8665w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range8550w8664w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9197w9393w9394w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9197w9393w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9329w9391w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9256w9475w9476w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9256w9475w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9358w9474w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9262w9483w9484w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9262w9483w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9361w9482w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9268w9491w9492w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9268w9491w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9364w9490w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9274w9499w9500w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9274w9499w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9367w9498w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9280w9507w9508w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9280w9507w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9370w9506w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9286w9515w9516w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9286w9515w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9373w9514w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9292w9523w9524w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9292w9523w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9376w9522w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9298w9531w9532w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9298w9531w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9379w9530w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9304w9539w9540w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9304w9539w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9382w9538w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9310w9547w9548w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9310w9547w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9385w9546w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9202w9403w9404w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9202w9403w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9331w9402w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9316w9555w9556w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9316w9555w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9388w9554w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9322w9563w9564w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9322w9563w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9167w9562w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9326w9571w9572w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9326w9571w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9171w9570w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9142w9579w9580w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9142w9579w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9173w9578w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9147w9587w9588w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9147w9587w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9175w9586w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9149w9595w9596w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9149w9595w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9177w9594w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9151w9603w9604w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9151w9603w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9179w9602w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9153w9611w9612w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9153w9611w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9181w9610w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9155w9619w9620w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9155w9619w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9183w9618w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9157w9627w9628w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9157w9627w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9185w9626w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9208w9411w9412w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9208w9411w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9334w9410w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9159w9635w9636w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9159w9635w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9187w9634w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9161w9643w9644w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9161w9643w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9189w9642w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9163w9651w9652w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9163w9651w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9191w9650w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9165w9659w9660w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9165w9659w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9193w9658w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9214w9419w9420w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9214w9419w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9337w9418w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9220w9427w9428w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9220w9427w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9340w9426w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9226w9435w9436w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9226w9435w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9343w9434w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9232w9443w9444w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9232w9443w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9346w9442w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9238w9451w9452w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9238w9451w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9349w9450w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9244w9459w9460w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9244w9459w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9352w9458w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9250w9467w9468w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range9250w9467w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range9355w9466w(0);
	wire_ccc_cordic_m_w10191w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10003w10190w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10129w10188w(0);
	wire_ccc_cordic_m_w10273w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10062w10272w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10158w10271w(0);
	wire_ccc_cordic_m_w10281w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10068w10280w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10161w10279w(0);
	wire_ccc_cordic_m_w10289w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10074w10288w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10164w10287w(0);
	wire_ccc_cordic_m_w10297w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10080w10296w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10167w10295w(0);
	wire_ccc_cordic_m_w10305w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10086w10304w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10170w10303w(0);
	wire_ccc_cordic_m_w10313w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10092w10312w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10173w10311w(0);
	wire_ccc_cordic_m_w10321w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10098w10320w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10176w10319w(0);
	wire_ccc_cordic_m_w10329w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10104w10328w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10179w10327w(0);
	wire_ccc_cordic_m_w10337w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10110w10336w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10182w10335w(0);
	wire_ccc_cordic_m_w10345w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10116w10344w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10185w10343w(0);
	wire_ccc_cordic_m_w10201w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10008w10200w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10131w10199w(0);
	wire_ccc_cordic_m_w10353w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10122w10352w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9971w10351w(0);
	wire_ccc_cordic_m_w10361w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10126w10360w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9975w10359w(0);
	wire_ccc_cordic_m_w10369w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9944w10368w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9977w10367w(0);
	wire_ccc_cordic_m_w10377w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9949w10376w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9979w10375w(0);
	wire_ccc_cordic_m_w10385w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9951w10384w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9981w10383w(0);
	wire_ccc_cordic_m_w10393w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9953w10392w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9983w10391w(0);
	wire_ccc_cordic_m_w10401w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9955w10400w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9985w10399w(0);
	wire_ccc_cordic_m_w10409w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9957w10408w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9987w10407w(0);
	wire_ccc_cordic_m_w10417w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9959w10416w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9989w10415w(0);
	wire_ccc_cordic_m_w10425w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9961w10424w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9991w10423w(0);
	wire_ccc_cordic_m_w10209w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10014w10208w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10134w10207w(0);
	wire_ccc_cordic_m_w10433w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9963w10432w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9993w10431w(0);
	wire_ccc_cordic_m_w10441w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9965w10440w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9995w10439w(0);
	wire_ccc_cordic_m_w10449w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9967w10448w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9997w10447w(0);
	wire_ccc_cordic_m_w10457w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9969w10456w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9999w10455w(0);
	wire_ccc_cordic_m_w10217w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10020w10216w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10137w10215w(0);
	wire_ccc_cordic_m_w10225w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10026w10224w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10140w10223w(0);
	wire_ccc_cordic_m_w10233w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10032w10232w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10143w10231w(0);
	wire_ccc_cordic_m_w10241w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10038w10240w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10146w10239w(0);
	wire_ccc_cordic_m_w10249w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10044w10248w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10149w10247w(0);
	wire_ccc_cordic_m_w10257w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10050w10256w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10152w10255w(0);
	wire_ccc_cordic_m_w10265w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range10056w10264w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range10155w10263w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range862w1148w1149w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range862w1148w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1054w1146w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range921w1230w1231w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range921w1230w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1083w1229w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range927w1238w1239w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range927w1238w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1086w1237w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range933w1246w1247w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range933w1246w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1089w1245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range939w1254w1255w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range939w1254w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1092w1253w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range945w1262w1263w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range945w1262w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1095w1261w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range951w1270w1271w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range951w1270w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1098w1269w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range957w1278w1279w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range957w1278w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1101w1277w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range963w1286w1287w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range963w1286w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1104w1285w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range969w1294w1295w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range969w1294w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1107w1293w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range975w1302w1303w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range975w1302w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1110w1301w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range867w1158w1159w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range867w1158w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1056w1157w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range981w1310w1311w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range981w1310w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1113w1309w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range987w1318w1319w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range987w1318w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1116w1317w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range993w1326w1327w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range993w1326w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1119w1325w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range999w1334w1335w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range999w1334w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1122w1333w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1005w1342w1343w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1005w1342w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1125w1341w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1011w1350w1351w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1011w1350w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1128w1349w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1017w1358w1359w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1017w1358w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1131w1357w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1023w1366w1367w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1023w1366w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1134w1365w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1029w1374w1375w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1029w1374w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1137w1373w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1035w1382w1383w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1035w1382w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1140w1381w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range873w1166w1167w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range873w1166w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1059w1165w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1041w1390w1391w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1041w1390w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1143w1389w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1047w1398w1399w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1047w1398w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range852w1397w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1051w1406w1407w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range1051w1406w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range856w1405w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range847w1414w1415w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range847w1414w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range858w1413w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range879w1174w1175w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range879w1174w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1062w1173w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range885w1182w1183w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range885w1182w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1065w1181w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range891w1190w1191w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range891w1190w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1068w1189w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range897w1198w1199w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range897w1198w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1071w1197w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range903w1206w1207w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range903w1206w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1074w1205w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range909w1214w1215w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range909w1214w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1077w1213w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range915w1222w1223w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range915w1222w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range1080w1221w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1718w1995w1996w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1718w1995w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1904w1993w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1777w2077w2078w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1777w2077w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1933w2076w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1783w2085w2086w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1783w2085w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1936w2084w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1789w2093w2094w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1789w2093w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1939w2092w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1795w2101w2102w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1795w2101w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1942w2100w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1801w2109w2110w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1801w2109w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1945w2108w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1807w2117w2118w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1807w2117w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1948w2116w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1813w2125w2126w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1813w2125w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1951w2124w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1819w2133w2134w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1819w2133w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1954w2132w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1825w2141w2142w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1825w2141w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1957w2140w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1831w2149w2150w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1831w2149w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1960w2148w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1723w2005w2006w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1723w2005w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1906w2004w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1837w2157w2158w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1837w2157w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1963w2156w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1843w2165w2166w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1843w2165w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1966w2164w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1849w2173w2174w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1849w2173w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1969w2172w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1855w2181w2182w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1855w2181w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1972w2180w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1861w2189w2190w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1861w2189w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1975w2188w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1867w2197w2198w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1867w2197w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1978w2196w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1873w2205w2206w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1873w2205w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1981w2204w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1879w2213w2214w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1879w2213w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1984w2212w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1885w2221w2222w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1885w2221w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1987w2220w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1891w2229w2230w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1891w2229w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1990w2228w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1729w2013w2014w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1729w2013w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1909w2012w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1897w2237w2238w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1897w2237w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1706w2236w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1901w2245w2246w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1901w2245w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1710w2244w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1699w2253w2254w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1699w2253w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1712w2252w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1704w2261w2262w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1704w2261w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1714w2260w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1735w2021w2022w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1735w2021w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1912w2020w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1741w2029w2030w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1741w2029w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1915w2028w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1747w2037w2038w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1747w2037w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1918w2036w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1753w2045w2046w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1753w2045w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1921w2044w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1759w2053w2054w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1759w2053w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1924w2052w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1765w2061w2062w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1765w2061w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1927w2060w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1771w2069w2070w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1771w2069w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1930w2068w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2569w2837w2838w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2569w2837w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2749w2835w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2628w2919w2920w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2628w2919w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2778w2918w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2634w2927w2928w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2634w2927w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2781w2926w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2640w2935w2936w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2640w2935w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2784w2934w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2646w2943w2944w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2646w2943w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2787w2942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2652w2951w2952w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2652w2951w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2790w2950w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2658w2959w2960w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2658w2959w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2793w2958w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2664w2967w2968w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2664w2967w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2796w2966w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2670w2975w2976w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2670w2975w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2799w2974w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2676w2983w2984w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2676w2983w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2802w2982w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2682w2991w2992w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2682w2991w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2805w2990w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2574w2847w2848w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2574w2847w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2751w2846w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2688w2999w3000w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2688w2999w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2808w2998w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2694w3007w3008w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2694w3007w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2811w3006w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2700w3015w3016w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2700w3015w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2814w3014w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2706w3023w3024w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2706w3023w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2817w3022w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2712w3031w3032w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2712w3031w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2820w3030w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2718w3039w3040w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2718w3039w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2823w3038w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2724w3047w3048w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2724w3047w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2826w3046w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2730w3055w3056w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2730w3055w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2829w3054w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2736w3063w3064w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2736w3063w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2832w3062w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2742w3071w3072w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2742w3071w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2555w3070w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2580w2855w2856w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2580w2855w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2754w2854w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2746w3079w3080w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2746w3079w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2559w3078w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2546w3087w3088w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2546w3087w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2561w3086w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2551w3095w3096w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2551w3095w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2563w3094w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2553w3103w3104w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2553w3103w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2565w3102w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2586w2863w2864w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2586w2863w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2757w2862w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2592w2871w2872w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2592w2871w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2760w2870w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2598w2879w2880w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2598w2879w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2763w2878w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2604w2887w2888w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2604w2887w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2766w2886w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2610w2895w2896w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2610w2895w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2769w2894w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2616w2903w2904w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2616w2903w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2772w2902w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2622w2911w2912w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2622w2911w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2775w2910w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3415w3674w3675w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3415w3674w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3589w3672w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3474w3756w3757w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3474w3756w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3618w3755w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3480w3764w3765w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3480w3764w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3621w3763w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3486w3772w3773w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3486w3772w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3624w3771w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3492w3780w3781w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3492w3780w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3627w3779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3498w3788w3789w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3498w3788w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3630w3787w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3504w3796w3797w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3504w3796w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3633w3795w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3510w3804w3805w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3510w3804w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3636w3803w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3516w3812w3813w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3516w3812w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3639w3811w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3522w3820w3821w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3522w3820w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3642w3819w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3528w3828w3829w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3528w3828w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3645w3827w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3420w3684w3685w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3420w3684w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3591w3683w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3534w3836w3837w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3534w3836w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3648w3835w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3540w3844w3845w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3540w3844w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3651w3843w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3546w3852w3853w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3546w3852w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3654w3851w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3552w3860w3861w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3552w3860w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3657w3859w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3558w3868w3869w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3558w3868w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3660w3867w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3564w3876w3877w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3564w3876w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3663w3875w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3570w3884w3885w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3570w3884w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3666w3883w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3576w3892w3893w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3576w3892w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3669w3891w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3582w3900w3901w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3582w3900w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3399w3899w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3586w3908w3909w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3586w3908w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3403w3907w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3426w3692w3693w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3426w3692w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3594w3691w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3388w3916w3917w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3388w3916w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3405w3915w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3393w3924w3925w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3393w3924w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3407w3923w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3395w3932w3933w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3395w3932w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3409w3931w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3397w3940w3941w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3397w3940w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3411w3939w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3432w3700w3701w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3432w3700w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3597w3699w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3438w3708w3709w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3438w3708w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3600w3707w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3444w3716w3717w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3444w3716w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3603w3715w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3450w3724w3725w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3450w3724w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3606w3723w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3456w3732w3733w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3456w3732w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3609w3731w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3462w3740w3741w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3462w3740w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3612w3739w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3468w3748w3749w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3468w3748w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3615w3747w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4256w4506w4507w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4256w4506w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4424w4504w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4315w4588w4589w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4315w4588w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4453w4587w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4321w4596w4597w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4321w4596w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4456w4595w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4327w4604w4605w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4327w4604w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4459w4603w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4333w4612w4613w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4333w4612w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4462w4611w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4339w4620w4621w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4339w4620w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4465w4619w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4345w4628w4629w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4345w4628w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4468w4627w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4351w4636w4637w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4351w4636w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4471w4635w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4357w4644w4645w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4357w4644w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4474w4643w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4363w4652w4653w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4363w4652w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4477w4651w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4369w4660w4661w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4369w4660w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4480w4659w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4261w4516w4517w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4261w4516w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4426w4515w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4375w4668w4669w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4375w4668w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4483w4667w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4381w4676w4677w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4381w4676w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4486w4675w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4387w4684w4685w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4387w4684w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4489w4683w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4393w4692w4693w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4393w4692w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4492w4691w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4399w4700w4701w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4399w4700w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4495w4699w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4405w4708w4709w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4405w4708w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4498w4707w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4411w4716w4717w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4411w4716w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4501w4715w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4417w4724w4725w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4417w4724w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4238w4723w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4421w4732w4733w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4421w4732w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4242w4731w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4225w4740w4741w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4225w4740w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4244w4739w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4267w4524w4525w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4267w4524w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4429w4523w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4230w4748w4749w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4230w4748w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4246w4747w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4232w4756w4757w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4232w4756w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4248w4755w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4234w4764w4765w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4234w4764w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4250w4763w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4236w4772w4773w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4236w4772w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4252w4771w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4273w4532w4533w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4273w4532w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4432w4531w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4279w4540w4541w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4279w4540w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4435w4539w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4285w4548w4549w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4285w4548w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4438w4547w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4291w4556w4557w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4291w4556w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4441w4555w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4297w4564w4565w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4297w4564w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4444w4563w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4303w4572w4573w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4303w4572w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4447w4571w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4309w4580w4581w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4309w4580w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4450w4579w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5092w5333w5334w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5092w5333w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5254w5331w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5151w5415w5416w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5151w5415w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5283w5414w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5157w5423w5424w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5157w5423w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5286w5422w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5163w5431w5432w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5163w5431w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5289w5430w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5169w5439w5440w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5169w5439w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5292w5438w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5175w5447w5448w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5175w5447w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5295w5446w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5181w5455w5456w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5181w5455w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5298w5454w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5187w5463w5464w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5187w5463w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5301w5462w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5193w5471w5472w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5193w5471w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5304w5470w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5199w5479w5480w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5199w5479w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5307w5478w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5205w5487w5488w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5205w5487w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5310w5486w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5097w5343w5344w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5097w5343w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5256w5342w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5211w5495w5496w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5211w5495w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5313w5494w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5217w5503w5504w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5217w5503w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5316w5502w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5223w5511w5512w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5223w5511w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5319w5510w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5229w5519w5520w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5229w5519w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5322w5518w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5235w5527w5528w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5235w5527w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5325w5526w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5241w5535w5536w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5241w5535w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5328w5534w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5247w5543w5544w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5247w5543w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5072w5542w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5251w5551w5552w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5251w5551w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5076w5550w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5057w5559w5560w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5057w5559w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5078w5558w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5062w5567w5568w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5062w5567w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5080w5566w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5103w5351w5352w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5103w5351w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5259w5350w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5064w5575w5576w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5064w5575w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5082w5574w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5066w5583w5584w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5066w5583w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5084w5582w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5068w5591w5592w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5068w5591w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5086w5590w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5070w5599w5600w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5070w5599w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5088w5598w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5109w5359w5360w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5109w5359w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5262w5358w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5115w5367w5368w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5115w5367w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5265w5366w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5121w5375w5376w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5121w5375w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5268w5374w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5127w5383w5384w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5127w5383w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5271w5382w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5133w5391w5392w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5133w5391w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5274w5390w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5139w5399w5400w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5139w5399w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5277w5398w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5145w5407w5408w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range5145w5407w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range5280w5406w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5923w6155w6156w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5923w6155w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6079w6153w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5982w6237w6238w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5982w6237w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6108w6236w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5988w6245w6246w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5988w6245w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6111w6244w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5994w6253w6254w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5994w6253w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6114w6252w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6000w6261w6262w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6000w6261w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6117w6260w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6006w6269w6270w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6006w6269w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6120w6268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6012w6277w6278w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6012w6277w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6123w6276w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6018w6285w6286w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6018w6285w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6126w6284w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6024w6293w6294w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6024w6293w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6129w6292w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6030w6301w6302w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6030w6301w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6132w6300w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6036w6309w6310w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6036w6309w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6135w6308w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5928w6165w6166w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5928w6165w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6081w6164w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6042w6317w6318w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6042w6317w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6138w6316w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6048w6325w6326w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6048w6325w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6141w6324w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6054w6333w6334w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6054w6333w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6144w6332w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6060w6341w6342w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6060w6341w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6147w6340w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6066w6349w6350w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6066w6349w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6150w6348w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6072w6357w6358w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6072w6357w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5901w6356w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6076w6365w6366w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range6076w6365w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5905w6364w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5884w6373w6374w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5884w6373w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5907w6372w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5889w6381w6382w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5889w6381w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5909w6380w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5891w6389w6390w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5891w6389w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5911w6388w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5934w6173w6174w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5934w6173w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6084w6172w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5893w6397w6398w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5893w6397w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5913w6396w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5895w6405w6406w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5895w6405w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5915w6404w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5897w6413w6414w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5897w6413w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5917w6412w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5899w6421w6422w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5899w6421w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5919w6420w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5940w6181w6182w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5940w6181w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6087w6180w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5946w6189w6190w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5946w6189w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6090w6188w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5952w6197w6198w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5952w6197w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6093w6196w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5958w6205w6206w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5958w6205w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6096w6204w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5964w6213w6214w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5964w6213w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6099w6212w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5970w6221w6222w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5970w6221w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6102w6220w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5976w6229w6230w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5976w6229w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range6105w6228w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6749w6972w6973w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6749w6972w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6899w6970w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6808w7054w7055w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6808w7054w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6928w7053w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6814w7062w7063w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6814w7062w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6931w7061w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6820w7070w7071w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6820w7070w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6934w7069w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6826w7078w7079w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6826w7078w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6937w7077w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6832w7086w7087w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6832w7086w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6940w7085w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6838w7094w7095w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6838w7094w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6943w7093w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6844w7102w7103w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6844w7102w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6946w7101w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6850w7110w7111w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6850w7110w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6949w7109w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6856w7118w7119w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6856w7118w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6952w7117w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6862w7126w7127w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6862w7126w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6955w7125w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6754w6982w6983w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6754w6982w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6901w6981w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6868w7134w7135w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6868w7134w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6958w7133w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6874w7142w7143w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6874w7142w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6961w7141w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6880w7150w7151w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6880w7150w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6964w7149w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6886w7158w7159w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6886w7158w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6967w7157w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6892w7166w7167w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6892w7166w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6725w7165w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6896w7174w7175w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6896w7174w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6729w7173w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6706w7182w7183w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6706w7182w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6731w7181w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6711w7190w7191w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6711w7190w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6733w7189w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6713w7198w7199w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6713w7198w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6735w7197w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6715w7206w7207w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6715w7206w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6737w7205w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6760w6990w6991w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6760w6990w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6904w6989w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6717w7214w7215w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6717w7214w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6739w7213w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6719w7222w7223w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6719w7222w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6741w7221w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6721w7230w7231w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6721w7230w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6743w7229w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6723w7238w7239w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6723w7238w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6745w7237w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6766w6998w6999w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6766w6998w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6907w6997w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6772w7006w7007w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6772w7006w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6910w7005w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6778w7014w7015w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6778w7014w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6913w7013w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6784w7022w7023w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6784w7022w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6916w7021w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6790w7030w7031w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6790w7030w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6919w7029w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6796w7038w7039w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6796w7038w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6922w7037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6802w7046w7047w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6802w7046w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6925w7045w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7572w7789w7790w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7572w7789w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7715w7788w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7631w7870w7871w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7631w7870w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7744w7869w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7637w7878w7879w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7637w7878w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7747w7877w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7643w7886w7887w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7643w7886w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7750w7885w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7649w7894w7895w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7649w7894w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7753w7893w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7655w7902w7903w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7655w7902w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7756w7901w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7661w7910w7911w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7661w7910w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7759w7909w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7667w7918w7919w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7667w7918w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7762w7917w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7673w7926w7927w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7673w7926w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7765w7925w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7679w7934w7935w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7679w7934w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7768w7933w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7685w7942w7943w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7685w7942w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7771w7941w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7577w7798w7799w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7577w7798w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7717w7797w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7691w7950w7951w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7691w7950w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7774w7949w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7697w7958w7959w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7697w7958w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7777w7957w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7703w7966w7967w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7703w7966w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7780w7965w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7709w7974w7975w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7709w7974w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7546w7973w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7712w7982w7983w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7712w7982w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7549w7981w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7526w7990w7991w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7526w7990w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7551w7989w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7529w7998w7999w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7529w7998w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7553w7997w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7531w8006w8007w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7531w8006w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7555w8005w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7533w8014w8015w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7533w8014w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7557w8013w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7535w8022w8023w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7535w8022w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7559w8021w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7583w7806w7807w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7583w7806w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7720w7805w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7537w8030w8031w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7537w8030w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7561w8029w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7539w8038w8039w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7539w8038w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7563w8037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7541w8046w8047w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7541w8046w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7565w8045w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7543w8054w8055w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7543w8054w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7567w8053w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7589w7814w7815w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7589w7814w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7723w7813w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7595w7822w7823w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7595w7822w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7726w7821w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7601w7830w7831w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7601w7830w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7729w7829w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7607w7838w7839w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7607w7838w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7732w7837w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7613w7846w7847w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7613w7846w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7735w7845w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7619w7854w7855w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7619w7854w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7738w7853w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7625w7862w7863w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7625w7862w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7741w7861w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8388w8596w8597w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8388w8596w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8525w8595w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8447w8677w8678w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8447w8677w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8554w8676w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8453w8685w8686w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8453w8685w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8557w8684w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8459w8693w8694w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8459w8693w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8560w8692w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8465w8701w8702w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8465w8701w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8563w8700w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8471w8709w8710w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8471w8709w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8566w8708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8477w8717w8718w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8477w8717w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8569w8716w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8483w8725w8726w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8483w8725w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8572w8724w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8489w8733w8734w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8489w8733w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8575w8732w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8495w8741w8742w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8495w8741w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8578w8740w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8501w8749w8750w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8501w8749w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8581w8748w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8393w8605w8606w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8393w8605w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8527w8604w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8507w8757w8758w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8507w8757w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8584w8756w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8513w8765w8766w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8513w8765w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8587w8764w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8519w8773w8774w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8519w8773w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8360w8772w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8522w8781w8782w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8522w8781w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8363w8780w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8338w8789w8790w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8338w8789w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8365w8788w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8341w8797w8798w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8341w8797w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8367w8796w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8343w8805w8806w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8343w8805w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8369w8804w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8345w8813w8814w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8345w8813w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8371w8812w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8347w8821w8822w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8347w8821w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8373w8820w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8349w8829w8830w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8349w8829w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8375w8828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8399w8613w8614w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8399w8613w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8530w8612w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8351w8837w8838w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8351w8837w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8377w8836w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8353w8845w8846w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8353w8845w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8379w8844w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8355w8853w8854w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8355w8853w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8381w8852w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8357w8861w8862w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8357w8861w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8383w8860w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8405w8621w8622w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8405w8621w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8533w8620w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8411w8629w8630w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8411w8629w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8536w8628w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8417w8637w8638w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8417w8637w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8539w8636w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8423w8645w8646w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8423w8645w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8542w8644w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8429w8653w8654w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8429w8653w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8545w8652w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8435w8661w8662w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8435w8661w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8548w8660w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8441w8669w8670w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range8441w8669w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range8551w8668w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9199w9398w9399w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9199w9398w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9330w9397w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9258w9479w9480w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9258w9479w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9359w9478w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9264w9487w9488w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9264w9487w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9362w9486w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9270w9495w9496w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9270w9495w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9365w9494w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9276w9503w9504w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9276w9503w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9368w9502w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9282w9511w9512w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9282w9511w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9371w9510w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9288w9519w9520w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9288w9519w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9374w9518w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9294w9527w9528w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9294w9527w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9377w9526w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9300w9535w9536w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9300w9535w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9380w9534w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9306w9543w9544w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9306w9543w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9383w9542w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9312w9551w9552w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9312w9551w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9386w9550w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9204w9407w9408w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9204w9407w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9332w9406w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9318w9559w9560w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9318w9559w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9389w9558w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9324w9567w9568w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9324w9567w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9169w9566w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9327w9575w9576w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9327w9575w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9172w9574w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9145w9583w9584w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9145w9583w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9174w9582w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9148w9591w9592w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9148w9591w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9176w9590w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9150w9599w9600w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9150w9599w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9178w9598w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9152w9607w9608w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9152w9607w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9180w9606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9154w9615w9616w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9154w9615w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9182w9614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9156w9623w9624w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9156w9623w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9184w9622w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9158w9631w9632w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9158w9631w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9186w9630w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9210w9415w9416w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9210w9415w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9335w9414w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9160w9639w9640w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9160w9639w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9188w9638w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9162w9647w9648w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9162w9647w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9190w9646w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9164w9655w9656w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9164w9655w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9192w9654w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9166w9663w9664w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9166w9663w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9194w9662w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9216w9423w9424w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9216w9423w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9338w9422w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9222w9431w9432w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9222w9431w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9341w9430w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9228w9439w9440w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9228w9439w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9344w9438w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9234w9447w9448w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9234w9447w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9347w9446w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9240w9455w9456w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9240w9455w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9350w9454w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9246w9463w9464w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9246w9463w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9353w9462w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9252w9471w9472w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range9252w9471w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range9356w9470w(0);
	wire_ccc_cordic_m_w10196w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10005w10195w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10130w10194w(0);
	wire_ccc_cordic_m_w10277w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10064w10276w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10159w10275w(0);
	wire_ccc_cordic_m_w10285w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10070w10284w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10162w10283w(0);
	wire_ccc_cordic_m_w10293w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10076w10292w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10165w10291w(0);
	wire_ccc_cordic_m_w10301w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10082w10300w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10168w10299w(0);
	wire_ccc_cordic_m_w10309w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10088w10308w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10171w10307w(0);
	wire_ccc_cordic_m_w10317w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10094w10316w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10174w10315w(0);
	wire_ccc_cordic_m_w10325w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10100w10324w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10177w10323w(0);
	wire_ccc_cordic_m_w10333w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10106w10332w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10180w10331w(0);
	wire_ccc_cordic_m_w10341w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10112w10340w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10183w10339w(0);
	wire_ccc_cordic_m_w10349w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10118w10348w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10186w10347w(0);
	wire_ccc_cordic_m_w10205w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10010w10204w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10132w10203w(0);
	wire_ccc_cordic_m_w10357w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10124w10356w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9973w10355w(0);
	wire_ccc_cordic_m_w10365w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10127w10364w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9976w10363w(0);
	wire_ccc_cordic_m_w10373w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9947w10372w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9978w10371w(0);
	wire_ccc_cordic_m_w10381w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9950w10380w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9980w10379w(0);
	wire_ccc_cordic_m_w10389w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9952w10388w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9982w10387w(0);
	wire_ccc_cordic_m_w10397w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9954w10396w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9984w10395w(0);
	wire_ccc_cordic_m_w10405w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9956w10404w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9986w10403w(0);
	wire_ccc_cordic_m_w10413w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9958w10412w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9988w10411w(0);
	wire_ccc_cordic_m_w10421w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9960w10420w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9990w10419w(0);
	wire_ccc_cordic_m_w10429w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9962w10428w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9992w10427w(0);
	wire_ccc_cordic_m_w10213w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10016w10212w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10135w10211w(0);
	wire_ccc_cordic_m_w10437w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9964w10436w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9994w10435w(0);
	wire_ccc_cordic_m_w10445w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9966w10444w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9996w10443w(0);
	wire_ccc_cordic_m_w10453w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9968w10452w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9998w10451w(0);
	wire_ccc_cordic_m_w10461w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9970w10460w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10000w10459w(0);
	wire_ccc_cordic_m_w10221w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10022w10220w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10138w10219w(0);
	wire_ccc_cordic_m_w10229w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10028w10228w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10141w10227w(0);
	wire_ccc_cordic_m_w10237w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10034w10236w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10144w10235w(0);
	wire_ccc_cordic_m_w10245w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10040w10244w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10147w10243w(0);
	wire_ccc_cordic_m_w10253w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10046w10252w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10150w10251w(0);
	wire_ccc_cordic_m_w10261w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10052w10260w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10153w10259w(0);
	wire_ccc_cordic_m_w10269w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range10058w10268w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range10156w10267w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range864w1153w1154w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range864w1153w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1055w1152w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range923w1234w1235w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range923w1234w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1084w1233w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range929w1242w1243w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range929w1242w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1087w1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range935w1250w1251w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range935w1250w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1090w1249w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range941w1258w1259w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range941w1258w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1093w1257w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range947w1266w1267w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range947w1266w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1096w1265w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range953w1274w1275w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range953w1274w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1099w1273w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range959w1282w1283w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range959w1282w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1102w1281w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range965w1290w1291w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range965w1290w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1105w1289w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range971w1298w1299w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range971w1298w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1108w1297w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range977w1306w1307w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range977w1306w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1111w1305w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range869w1162w1163w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range869w1162w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1057w1161w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range983w1314w1315w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range983w1314w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1114w1313w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range989w1322w1323w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range989w1322w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1117w1321w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range995w1330w1331w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range995w1330w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1120w1329w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1001w1338w1339w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1001w1338w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1123w1337w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1007w1346w1347w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1007w1346w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1126w1345w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1013w1354w1355w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1013w1354w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1129w1353w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1019w1362w1363w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1019w1362w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1132w1361w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1025w1370w1371w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1025w1370w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1135w1369w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1031w1378w1379w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1031w1378w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1138w1377w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1037w1386w1387w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1037w1386w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1141w1385w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range875w1170w1171w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range875w1170w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1060w1169w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1043w1394w1395w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1043w1394w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1144w1393w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1049w1402w1403w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1049w1402w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range854w1401w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1052w1410w1411w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range1052w1410w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range857w1409w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range850w1418w1419w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range850w1418w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range859w1417w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range881w1178w1179w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range881w1178w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1063w1177w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range887w1186w1187w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range887w1186w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1066w1185w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range893w1194w1195w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range893w1194w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1069w1193w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range899w1202w1203w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range899w1202w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1072w1201w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range905w1210w1211w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range905w1210w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1075w1209w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range911w1218w1219w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range911w1218w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1078w1217w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range917w1226w1227w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range917w1226w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range1081w1225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1720w2000w2001w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1720w2000w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1905w1999w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1779w2081w2082w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1779w2081w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1934w2080w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1785w2089w2090w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1785w2089w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1937w2088w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1791w2097w2098w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1791w2097w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1940w2096w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1797w2105w2106w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1797w2105w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1943w2104w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1803w2113w2114w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1803w2113w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1946w2112w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1809w2121w2122w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1809w2121w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1949w2120w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1815w2129w2130w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1815w2129w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1952w2128w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1821w2137w2138w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1821w2137w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1955w2136w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1827w2145w2146w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1827w2145w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1958w2144w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1833w2153w2154w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1833w2153w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1961w2152w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1725w2009w2010w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1725w2009w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1907w2008w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1839w2161w2162w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1839w2161w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1964w2160w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1845w2169w2170w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1845w2169w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1967w2168w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1851w2177w2178w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1851w2177w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1970w2176w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1857w2185w2186w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1857w2185w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1973w2184w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1863w2193w2194w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1863w2193w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1976w2192w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1869w2201w2202w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1869w2201w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1979w2200w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1875w2209w2210w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1875w2209w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1982w2208w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1881w2217w2218w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1881w2217w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1985w2216w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1887w2225w2226w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1887w2225w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1988w2224w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1893w2233w2234w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1893w2233w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1991w2232w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1731w2017w2018w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1731w2017w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1910w2016w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1899w2241w2242w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1899w2241w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1708w2240w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1902w2249w2250w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1902w2249w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1711w2248w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1702w2257w2258w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1702w2257w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1713w2256w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1705w2265w2266w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1705w2265w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1715w2264w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1737w2025w2026w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1737w2025w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1913w2024w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1743w2033w2034w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1743w2033w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1916w2032w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1749w2041w2042w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1749w2041w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1919w2040w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1755w2049w2050w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1755w2049w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1922w2048w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1761w2057w2058w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1761w2057w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1925w2056w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1767w2065w2066w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1767w2065w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1928w2064w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1773w2073w2074w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1773w2073w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1931w2072w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2571w2842w2843w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2571w2842w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2750w2841w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2630w2923w2924w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2630w2923w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2779w2922w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2636w2931w2932w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2636w2931w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2782w2930w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2642w2939w2940w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2642w2939w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2785w2938w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2648w2947w2948w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2648w2947w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2788w2946w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2654w2955w2956w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2654w2955w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2791w2954w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2660w2963w2964w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2660w2963w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2794w2962w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2666w2971w2972w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2666w2971w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2797w2970w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2672w2979w2980w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2672w2979w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2800w2978w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2678w2987w2988w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2678w2987w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2803w2986w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2684w2995w2996w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2684w2995w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2806w2994w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2576w2851w2852w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2576w2851w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2752w2850w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2690w3003w3004w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2690w3003w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2809w3002w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2696w3011w3012w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2696w3011w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2812w3010w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2702w3019w3020w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2702w3019w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2815w3018w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2708w3027w3028w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2708w3027w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2818w3026w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2714w3035w3036w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2714w3035w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2821w3034w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2720w3043w3044w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2720w3043w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2824w3042w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2726w3051w3052w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2726w3051w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2827w3050w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2732w3059w3060w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2732w3059w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2830w3058w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2738w3067w3068w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2738w3067w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2833w3066w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2744w3075w3076w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2744w3075w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2557w3074w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2582w2859w2860w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2582w2859w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2755w2858w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2747w3083w3084w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2747w3083w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2560w3082w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2549w3091w3092w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2549w3091w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2562w3090w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2552w3099w3100w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2552w3099w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2564w3098w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2554w3107w3108w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2554w3107w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2566w3106w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2588w2867w2868w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2588w2867w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2758w2866w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2594w2875w2876w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2594w2875w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2761w2874w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2600w2883w2884w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2600w2883w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2764w2882w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2606w2891w2892w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2606w2891w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2767w2890w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2612w2899w2900w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2612w2899w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2770w2898w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2618w2907w2908w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2618w2907w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2773w2906w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2624w2915w2916w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2624w2915w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2776w2914w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3417w3679w3680w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3417w3679w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3590w3678w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3476w3760w3761w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3476w3760w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3619w3759w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3482w3768w3769w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3482w3768w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3622w3767w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3488w3776w3777w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3488w3776w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3625w3775w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3494w3784w3785w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3494w3784w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3628w3783w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3500w3792w3793w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3500w3792w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3631w3791w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3506w3800w3801w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3506w3800w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3634w3799w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3512w3808w3809w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3512w3808w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3637w3807w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3518w3816w3817w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3518w3816w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3640w3815w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3524w3824w3825w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3524w3824w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3643w3823w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3530w3832w3833w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3530w3832w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3646w3831w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3422w3688w3689w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3422w3688w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3592w3687w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3536w3840w3841w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3536w3840w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3649w3839w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3542w3848w3849w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3542w3848w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3652w3847w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3548w3856w3857w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3548w3856w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3655w3855w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3554w3864w3865w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3554w3864w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3658w3863w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3560w3872w3873w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3560w3872w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3661w3871w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3566w3880w3881w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3566w3880w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3664w3879w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3572w3888w3889w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3572w3888w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3667w3887w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3578w3896w3897w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3578w3896w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3670w3895w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3584w3904w3905w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3584w3904w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3401w3903w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3587w3912w3913w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3587w3912w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3404w3911w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3428w3696w3697w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3428w3696w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3595w3695w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3391w3920w3921w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3391w3920w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3406w3919w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3394w3928w3929w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3394w3928w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3408w3927w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3396w3936w3937w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3396w3936w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3410w3935w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3398w3944w3945w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3398w3944w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3412w3943w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3434w3704w3705w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3434w3704w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3598w3703w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3440w3712w3713w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3440w3712w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3601w3711w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3446w3720w3721w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3446w3720w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3604w3719w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3452w3728w3729w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3452w3728w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3607w3727w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3458w3736w3737w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3458w3736w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3610w3735w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3464w3744w3745w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3464w3744w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3613w3743w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3470w3752w3753w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3470w3752w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3616w3751w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4258w4511w4512w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4258w4511w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4425w4510w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4317w4592w4593w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4317w4592w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4454w4591w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4323w4600w4601w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4323w4600w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4457w4599w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4329w4608w4609w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4329w4608w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4460w4607w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4335w4616w4617w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4335w4616w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4463w4615w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4341w4624w4625w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4341w4624w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4466w4623w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4347w4632w4633w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4347w4632w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4469w4631w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4353w4640w4641w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4353w4640w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4472w4639w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4359w4648w4649w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4359w4648w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4475w4647w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4365w4656w4657w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4365w4656w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4478w4655w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4371w4664w4665w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4371w4664w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4481w4663w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4263w4520w4521w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4263w4520w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4427w4519w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4377w4672w4673w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4377w4672w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4484w4671w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4383w4680w4681w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4383w4680w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4487w4679w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4389w4688w4689w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4389w4688w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4490w4687w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4395w4696w4697w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4395w4696w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4493w4695w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4401w4704w4705w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4401w4704w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4496w4703w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4407w4712w4713w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4407w4712w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4499w4711w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4413w4720w4721w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4413w4720w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4502w4719w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4419w4728w4729w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4419w4728w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4240w4727w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4422w4736w4737w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4422w4736w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4243w4735w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4228w4744w4745w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4228w4744w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4245w4743w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4269w4528w4529w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4269w4528w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4430w4527w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4231w4752w4753w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4231w4752w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4247w4751w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4233w4760w4761w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4233w4760w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4249w4759w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4235w4768w4769w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4235w4768w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4251w4767w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4237w4776w4777w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4237w4776w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4253w4775w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4275w4536w4537w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4275w4536w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4433w4535w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4281w4544w4545w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4281w4544w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4436w4543w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4287w4552w4553w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4287w4552w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4439w4551w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4293w4560w4561w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4293w4560w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4442w4559w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4299w4568w4569w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4299w4568w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4445w4567w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4305w4576w4577w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4305w4576w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4448w4575w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4311w4584w4585w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4311w4584w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4451w4583w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5094w5338w5339w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5094w5338w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5255w5337w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5153w5419w5420w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5153w5419w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5284w5418w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5159w5427w5428w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5159w5427w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5287w5426w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5165w5435w5436w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5165w5435w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5290w5434w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5171w5443w5444w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5171w5443w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5293w5442w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5177w5451w5452w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5177w5451w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5296w5450w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5183w5459w5460w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5183w5459w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5299w5458w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5189w5467w5468w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5189w5467w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5302w5466w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5195w5475w5476w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5195w5475w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5305w5474w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5201w5483w5484w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5201w5483w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5308w5482w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5207w5491w5492w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5207w5491w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5311w5490w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5099w5347w5348w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5099w5347w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5257w5346w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5213w5499w5500w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5213w5499w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5314w5498w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5219w5507w5508w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5219w5507w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5317w5506w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5225w5515w5516w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5225w5515w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5320w5514w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5231w5523w5524w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5231w5523w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5323w5522w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5237w5531w5532w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5237w5531w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5326w5530w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5243w5539w5540w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5243w5539w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5329w5538w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5249w5547w5548w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5249w5547w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5074w5546w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5252w5555w5556w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5252w5555w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5077w5554w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5060w5563w5564w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5060w5563w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5079w5562w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5063w5571w5572w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5063w5571w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5081w5570w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5105w5355w5356w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5105w5355w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5260w5354w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5065w5579w5580w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5065w5579w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5083w5578w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5067w5587w5588w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5067w5587w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5085w5586w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5069w5595w5596w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5069w5595w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5087w5594w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5071w5603w5604w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5071w5603w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5089w5602w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5111w5363w5364w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5111w5363w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5263w5362w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5117w5371w5372w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5117w5371w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5266w5370w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5123w5379w5380w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5123w5379w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5269w5378w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5129w5387w5388w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5129w5387w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5272w5386w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5135w5395w5396w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5135w5395w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5275w5394w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5141w5403w5404w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5141w5403w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5278w5402w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5147w5411w5412w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range5147w5411w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range5281w5410w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5925w6160w6161w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5925w6160w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6080w6159w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5984w6241w6242w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5984w6241w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6109w6240w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5990w6249w6250w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5990w6249w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6112w6248w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5996w6257w6258w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5996w6257w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6115w6256w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6002w6265w6266w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6002w6265w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6118w6264w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6008w6273w6274w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6008w6273w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6121w6272w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6014w6281w6282w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6014w6281w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6124w6280w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6020w6289w6290w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6020w6289w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6127w6288w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6026w6297w6298w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6026w6297w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6130w6296w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6032w6305w6306w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6032w6305w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6133w6304w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6038w6313w6314w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6038w6313w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6136w6312w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5930w6169w6170w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5930w6169w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6082w6168w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6044w6321w6322w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6044w6321w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6139w6320w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6050w6329w6330w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6050w6329w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6142w6328w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6056w6337w6338w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6056w6337w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6145w6336w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6062w6345w6346w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6062w6345w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6148w6344w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6068w6353w6354w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6068w6353w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6151w6352w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6074w6361w6362w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6074w6361w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5903w6360w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6077w6369w6370w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range6077w6369w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5906w6368w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5887w6377w6378w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5887w6377w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5908w6376w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5890w6385w6386w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5890w6385w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5910w6384w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5892w6393w6394w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5892w6393w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5912w6392w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5936w6177w6178w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5936w6177w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6085w6176w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5894w6401w6402w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5894w6401w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5914w6400w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5896w6409w6410w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5896w6409w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5916w6408w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5898w6417w6418w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5898w6417w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5918w6416w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5900w6425w6426w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5900w6425w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5920w6424w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5942w6185w6186w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5942w6185w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6088w6184w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5948w6193w6194w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5948w6193w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6091w6192w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5954w6201w6202w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5954w6201w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6094w6200w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5960w6209w6210w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5960w6209w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6097w6208w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5966w6217w6218w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5966w6217w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6100w6216w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5972w6225w6226w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5972w6225w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6103w6224w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5978w6233w6234w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5978w6233w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range6106w6232w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6751w6977w6978w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6751w6977w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6900w6976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6810w7058w7059w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6810w7058w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6929w7057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6816w7066w7067w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6816w7066w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6932w7065w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6822w7074w7075w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6822w7074w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6935w7073w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6828w7082w7083w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6828w7082w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6938w7081w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6834w7090w7091w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6834w7090w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6941w7089w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6840w7098w7099w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6840w7098w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6944w7097w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6846w7106w7107w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6846w7106w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6947w7105w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6852w7114w7115w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6852w7114w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6950w7113w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6858w7122w7123w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6858w7122w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6953w7121w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6864w7130w7131w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6864w7130w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6956w7129w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6756w6986w6987w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6756w6986w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6902w6985w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6870w7138w7139w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6870w7138w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6959w7137w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6876w7146w7147w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6876w7146w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6962w7145w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6882w7154w7155w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6882w7154w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6965w7153w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6888w7162w7163w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6888w7162w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6968w7161w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6894w7170w7171w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6894w7170w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6727w7169w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6897w7178w7179w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6897w7178w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6730w7177w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6709w7186w7187w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6709w7186w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6732w7185w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6712w7194w7195w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6712w7194w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6734w7193w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6714w7202w7203w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6714w7202w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6736w7201w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6716w7210w7211w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6716w7210w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6738w7209w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6762w6994w6995w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6762w6994w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6905w6993w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6718w7218w7219w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6718w7218w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6740w7217w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6720w7226w7227w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6720w7226w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6742w7225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6722w7234w7235w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6722w7234w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6744w7233w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6724w7242w7243w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6724w7242w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6746w7241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6768w7002w7003w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6768w7002w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6908w7001w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6774w7010w7011w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6774w7010w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6911w7009w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6780w7018w7019w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6780w7018w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6914w7017w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6786w7026w7027w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6786w7026w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6917w7025w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6792w7034w7035w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6792w7034w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6920w7033w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6798w7042w7043w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6798w7042w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6923w7041w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6804w7050w7051w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6804w7050w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6926w7049w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8871w8872w8873w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8871w8872w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8952w8953w8954w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8952w8953w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8960w8961w8962w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8960w8961w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8968w8969w8970w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8968w8969w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8976w8977w8978w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8976w8977w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8984w8985w8986w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8984w8985w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8992w8993w8994w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8992w8993w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9000w9001w9002w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9000w9001w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9008w9009w9010w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9008w9009w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9016w9017w9018w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9016w9017w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9024w9025w9026w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9024w9025w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8880w8881w8882w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8880w8881w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9032w9033w9034w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9032w9033w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9040w9041w9042w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9040w9041w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9048w9049w9050w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9048w9049w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9056w9057w9058w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9056w9057w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9064w9065w9066w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9064w9065w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9072w9073w9074w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9072w9073w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9080w9081w9082w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9080w9081w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9088w9089w9090w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9088w9089w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9096w9097w9098w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9096w9097w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9104w9105w9106w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9104w9105w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8888w8889w8890w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8888w8889w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9112w9113w9114w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9112w9113w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9120w9121w9122w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9120w9121w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9128w9129w9130w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9128w9129w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9136w9137w9138w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range9136w9137w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8896w8897w8898w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8896w8897w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8904w8905w8906w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8904w8905w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8912w8913w8914w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8912w8913w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8920w8921w8922w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8920w8921w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8928w8929w8930w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8928w8929w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8936w8937w8938w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8936w8937w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8944w8945w8946w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8944w8945w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9673w9674w9675w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9673w9674w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9754w9755w9756w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9754w9755w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9762w9763w9764w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9762w9763w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9770w9771w9772w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9770w9771w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9778w9779w9780w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9778w9779w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9786w9787w9788w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9786w9787w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9794w9795w9796w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9794w9795w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9802w9803w9804w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9802w9803w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9810w9811w9812w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9810w9811w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9818w9819w9820w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9818w9819w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9826w9827w9828w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9826w9827w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9682w9683w9684w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9682w9683w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9834w9835w9836w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9834w9835w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9842w9843w9844w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9842w9843w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9850w9851w9852w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9850w9851w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9858w9859w9860w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9858w9859w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9866w9867w9868w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9866w9867w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9874w9875w9876w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9874w9875w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9882w9883w9884w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9882w9883w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9890w9891w9892w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9890w9891w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9898w9899w9900w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9898w9899w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9906w9907w9908w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9906w9907w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9690w9691w9692w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9690w9691w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9914w9915w9916w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9914w9915w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9922w9923w9924w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9922w9923w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9930w9931w9932w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9930w9931w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9938w9939w9940w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9938w9939w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9698w9699w9700w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9698w9699w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9706w9707w9708w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9706w9707w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9714w9715w9716w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9714w9715w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9722w9723w9724w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9722w9723w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9730w9731w9732w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9730w9731w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9738w9739w9740w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9738w9739w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9746w9747w9748w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9746w9747w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10470w10471w10472w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10470w10471w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10551w10552w10553w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10551w10552w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10559w10560w10561w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10559w10560w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10567w10568w10569w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10567w10568w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10575w10576w10577w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10575w10576w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10583w10584w10585w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10583w10584w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10591w10592w10593w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10591w10592w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10599w10600w10601w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10599w10600w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10607w10608w10609w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10607w10608w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10615w10616w10617w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10615w10616w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10623w10624w10625w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10623w10624w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10479w10480w10481w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10479w10480w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10631w10632w10633w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10631w10632w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10639w10640w10641w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10639w10640w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10647w10648w10649w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10647w10648w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10655w10656w10657w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10655w10656w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10663w10664w10665w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10663w10664w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10671w10672w10673w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10671w10672w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10679w10680w10681w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10679w10680w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10687w10688w10689w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10687w10688w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10695w10696w10697w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10695w10696w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10703w10704w10705w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10703w10704w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10487w10488w10489w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10487w10488w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10711w10712w10713w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10711w10712w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10719w10720w10721w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10719w10720w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10727w10728w10729w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10727w10728w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10735w10736w10737w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10735w10736w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10495w10496w10497w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10495w10496w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10503w10504w10505w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10503w10504w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10511w10512w10513w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10511w10512w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10519w10520w10521w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10519w10520w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10527w10528w10529w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10527w10528w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10535w10536w10537w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10535w10536w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10543w10544w10545w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range10543w10544w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1428w1429w1430w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1428w1429w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1509w1510w1511w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1509w1510w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1517w1518w1519w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1517w1518w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1525w1526w1527w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1525w1526w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1533w1534w1535w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1533w1534w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1541w1542w1543w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1541w1542w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1549w1550w1551w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1549w1550w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1557w1558w1559w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1557w1558w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1565w1566w1567w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1565w1566w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1573w1574w1575w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1573w1574w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1581w1582w1583w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1581w1582w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1437w1438w1439w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1437w1438w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1589w1590w1591w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1589w1590w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1597w1598w1599w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1597w1598w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1605w1606w1607w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1605w1606w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1613w1614w1615w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1613w1614w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1621w1622w1623w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1621w1622w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1629w1630w1631w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1629w1630w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1637w1638w1639w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1637w1638w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1645w1646w1647w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1645w1646w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1653w1654w1655w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1653w1654w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1661w1662w1663w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1661w1662w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1445w1446w1447w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1445w1446w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1669w1670w1671w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1669w1670w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1677w1678w1679w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1677w1678w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1685w1686w1687w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1685w1686w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1693w1694w1695w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1693w1694w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1453w1454w1455w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1453w1454w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1461w1462w1463w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1461w1462w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1469w1470w1471w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1469w1470w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1477w1478w1479w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1477w1478w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1485w1486w1487w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1485w1486w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1493w1494w1495w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1493w1494w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1501w1502w1503w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1501w1502w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2275w2276w2277w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2275w2276w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2356w2357w2358w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2356w2357w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2364w2365w2366w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2364w2365w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2372w2373w2374w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2372w2373w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2380w2381w2382w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2380w2381w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2388w2389w2390w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2388w2389w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2396w2397w2398w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2396w2397w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2404w2405w2406w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2404w2405w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2412w2413w2414w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2412w2413w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2420w2421w2422w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2420w2421w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2428w2429w2430w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2428w2429w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2284w2285w2286w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2284w2285w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2436w2437w2438w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2436w2437w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2444w2445w2446w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2444w2445w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2452w2453w2454w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2452w2453w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2460w2461w2462w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2460w2461w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2468w2469w2470w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2468w2469w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2476w2477w2478w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2476w2477w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2484w2485w2486w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2484w2485w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2492w2493w2494w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2492w2493w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2500w2501w2502w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2500w2501w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2508w2509w2510w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2508w2509w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2292w2293w2294w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2292w2293w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2516w2517w2518w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2516w2517w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2524w2525w2526w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2524w2525w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2532w2533w2534w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2532w2533w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2540w2541w2542w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2540w2541w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2300w2301w2302w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2300w2301w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2308w2309w2310w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2308w2309w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2316w2317w2318w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2316w2317w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2324w2325w2326w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2324w2325w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2332w2333w2334w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2332w2333w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2340w2341w2342w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2340w2341w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2348w2349w2350w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2348w2349w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3117w3118w3119w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3117w3118w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3198w3199w3200w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3198w3199w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3206w3207w3208w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3206w3207w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3214w3215w3216w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3214w3215w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3222w3223w3224w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3222w3223w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3230w3231w3232w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3230w3231w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3238w3239w3240w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3238w3239w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3246w3247w3248w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3246w3247w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3254w3255w3256w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3254w3255w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3262w3263w3264w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3262w3263w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3270w3271w3272w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3270w3271w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3126w3127w3128w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3126w3127w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3278w3279w3280w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3278w3279w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3286w3287w3288w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3286w3287w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3294w3295w3296w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3294w3295w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3302w3303w3304w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3302w3303w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3310w3311w3312w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3310w3311w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3318w3319w3320w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3318w3319w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3326w3327w3328w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3326w3327w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3334w3335w3336w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3334w3335w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3342w3343w3344w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3342w3343w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3350w3351w3352w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3350w3351w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3134w3135w3136w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3134w3135w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3358w3359w3360w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3358w3359w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3366w3367w3368w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3366w3367w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3374w3375w3376w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3374w3375w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3382w3383w3384w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3382w3383w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3142w3143w3144w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3142w3143w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3150w3151w3152w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3150w3151w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3158w3159w3160w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3158w3159w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3166w3167w3168w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3166w3167w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3174w3175w3176w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3174w3175w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3182w3183w3184w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3182w3183w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3190w3191w3192w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3190w3191w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3954w3955w3956w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3954w3955w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4035w4036w4037w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4035w4036w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4043w4044w4045w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4043w4044w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4051w4052w4053w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4051w4052w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4059w4060w4061w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4059w4060w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4067w4068w4069w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4067w4068w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4075w4076w4077w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4075w4076w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4083w4084w4085w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4083w4084w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4091w4092w4093w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4091w4092w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4099w4100w4101w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4099w4100w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4107w4108w4109w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4107w4108w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3963w3964w3965w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3963w3964w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4115w4116w4117w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4115w4116w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4123w4124w4125w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4123w4124w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4131w4132w4133w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4131w4132w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4139w4140w4141w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4139w4140w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4147w4148w4149w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4147w4148w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4155w4156w4157w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4155w4156w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4163w4164w4165w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4163w4164w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4171w4172w4173w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4171w4172w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4179w4180w4181w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4179w4180w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4187w4188w4189w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4187w4188w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3971w3972w3973w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3971w3972w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4195w4196w4197w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4195w4196w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4203w4204w4205w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4203w4204w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4211w4212w4213w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4211w4212w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4219w4220w4221w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4219w4220w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3979w3980w3981w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3979w3980w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3987w3988w3989w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3987w3988w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3995w3996w3997w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3995w3996w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4003w4004w4005w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4003w4004w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4011w4012w4013w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4011w4012w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4019w4020w4021w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4019w4020w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4027w4028w4029w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range4027w4028w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4786w4787w4788w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4786w4787w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4867w4868w4869w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4867w4868w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4875w4876w4877w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4875w4876w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4883w4884w4885w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4883w4884w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4891w4892w4893w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4891w4892w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4899w4900w4901w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4899w4900w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4907w4908w4909w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4907w4908w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4915w4916w4917w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4915w4916w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4923w4924w4925w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4923w4924w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4931w4932w4933w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4931w4932w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4939w4940w4941w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4939w4940w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4795w4796w4797w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4795w4796w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4947w4948w4949w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4947w4948w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4955w4956w4957w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4955w4956w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4963w4964w4965w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4963w4964w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4971w4972w4973w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4971w4972w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4979w4980w4981w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4979w4980w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4987w4988w4989w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4987w4988w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4995w4996w4997w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4995w4996w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5003w5004w5005w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5003w5004w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5011w5012w5013w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5011w5012w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5019w5020w5021w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5019w5020w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4803w4804w4805w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4803w4804w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5027w5028w5029w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5027w5028w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5035w5036w5037w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5035w5036w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5043w5044w5045w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5043w5044w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5051w5052w5053w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range5051w5052w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4811w4812w4813w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4811w4812w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4819w4820w4821w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4819w4820w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4827w4828w4829w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4827w4828w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4835w4836w4837w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4835w4836w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4843w4844w4845w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4843w4844w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4851w4852w4853w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4851w4852w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4859w4860w4861w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4859w4860w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5613w5614w5615w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5613w5614w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5694w5695w5696w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5694w5695w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5702w5703w5704w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5702w5703w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5710w5711w5712w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5710w5711w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5718w5719w5720w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5718w5719w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5726w5727w5728w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5726w5727w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5734w5735w5736w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5734w5735w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5742w5743w5744w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5742w5743w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5750w5751w5752w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5750w5751w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5758w5759w5760w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5758w5759w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5766w5767w5768w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5766w5767w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5622w5623w5624w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5622w5623w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5774w5775w5776w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5774w5775w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5782w5783w5784w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5782w5783w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5790w5791w5792w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5790w5791w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5798w5799w5800w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5798w5799w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5806w5807w5808w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5806w5807w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5814w5815w5816w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5814w5815w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5822w5823w5824w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5822w5823w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5830w5831w5832w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5830w5831w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5838w5839w5840w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5838w5839w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5846w5847w5848w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5846w5847w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5630w5631w5632w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5630w5631w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5854w5855w5856w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5854w5855w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5862w5863w5864w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5862w5863w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5870w5871w5872w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5870w5871w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5878w5879w5880w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5878w5879w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5638w5639w5640w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5638w5639w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5646w5647w5648w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5646w5647w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5654w5655w5656w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5654w5655w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5662w5663w5664w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5662w5663w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5670w5671w5672w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5670w5671w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5678w5679w5680w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5678w5679w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5686w5687w5688w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5686w5687w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6435w6436w6437w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6435w6436w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6516w6517w6518w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6516w6517w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6524w6525w6526w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6524w6525w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6532w6533w6534w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6532w6533w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6540w6541w6542w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6540w6541w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6548w6549w6550w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6548w6549w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6556w6557w6558w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6556w6557w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6564w6565w6566w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6564w6565w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6572w6573w6574w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6572w6573w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6580w6581w6582w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6580w6581w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6588w6589w6590w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6588w6589w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6444w6445w6446w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6444w6445w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6596w6597w6598w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6596w6597w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6604w6605w6606w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6604w6605w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6612w6613w6614w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6612w6613w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6620w6621w6622w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6620w6621w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6628w6629w6630w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6628w6629w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6636w6637w6638w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6636w6637w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6644w6645w6646w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6644w6645w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6652w6653w6654w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6652w6653w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6660w6661w6662w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6660w6661w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6668w6669w6670w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6668w6669w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6452w6453w6454w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6452w6453w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6676w6677w6678w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6676w6677w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6684w6685w6686w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6684w6685w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6692w6693w6694w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6692w6693w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6700w6701w6702w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6700w6701w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6460w6461w6462w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6460w6461w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6468w6469w6470w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6468w6469w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6476w6477w6478w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6476w6477w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6484w6485w6486w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6484w6485w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6492w6493w6494w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6492w6493w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6500w6501w6502w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6500w6501w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6508w6509w6510w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6508w6509w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7252w7253w7254w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7252w7253w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7333w7334w7335w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7333w7334w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7341w7342w7343w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7341w7342w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7349w7350w7351w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7349w7350w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7357w7358w7359w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7357w7358w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7365w7366w7367w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7365w7366w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7373w7374w7375w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7373w7374w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7381w7382w7383w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7381w7382w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7389w7390w7391w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7389w7390w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7397w7398w7399w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7397w7398w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7405w7406w7407w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7405w7406w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7261w7262w7263w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7261w7262w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7413w7414w7415w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7413w7414w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7421w7422w7423w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7421w7422w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7429w7430w7431w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7429w7430w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7437w7438w7439w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7437w7438w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7445w7446w7447w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7445w7446w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7453w7454w7455w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7453w7454w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7461w7462w7463w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7461w7462w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7469w7470w7471w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7469w7470w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7477w7478w7479w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7477w7478w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7485w7486w7487w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7485w7486w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7269w7270w7271w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7269w7270w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7493w7494w7495w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7493w7494w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7501w7502w7503w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7501w7502w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7509w7510w7511w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7509w7510w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7517w7518w7519w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7517w7518w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7277w7278w7279w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7277w7278w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7285w7286w7287w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7285w7286w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7293w7294w7295w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7293w7294w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7301w7302w7303w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7301w7302w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7309w7310w7311w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7309w7310w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7317w7318w7319w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7317w7318w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7325w7326w7327w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range7325w7326w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8064w8065w8066w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8064w8065w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8145w8146w8147w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8145w8146w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8153w8154w8155w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8153w8154w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8161w8162w8163w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8161w8162w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8169w8170w8171w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8169w8170w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8177w8178w8179w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8177w8178w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8185w8186w8187w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8185w8186w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8193w8194w8195w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8193w8194w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8201w8202w8203w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8201w8202w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8209w8210w8211w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8209w8210w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8217w8218w8219w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8217w8218w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8073w8074w8075w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8073w8074w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8225w8226w8227w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8225w8226w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8233w8234w8235w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8233w8234w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8241w8242w8243w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8241w8242w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8249w8250w8251w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8249w8250w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8257w8258w8259w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8257w8258w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8265w8266w8267w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8265w8266w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8273w8274w8275w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8273w8274w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8281w8282w8283w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8281w8282w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8289w8290w8291w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8289w8290w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8297w8298w8299w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8297w8298w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8081w8082w8083w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8081w8082w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8305w8306w8307w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8305w8306w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8313w8314w8315w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8313w8314w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8321w8322w8323w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8321w8322w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8329w8330w8331w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8329w8330w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8089w8090w8091w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8089w8090w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8097w8098w8099w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8097w8098w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8105w8106w8107w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8105w8106w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8113w8114w8115w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8113w8114w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8121w8122w8123w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8121w8122w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8129w8130w8131w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8129w8130w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8137w8138w8139w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range8137w8138w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	loop31 : FOR i IN 0 TO 33 GENERATE 
		wire_ccc_cordic_m_w_lg_estimate_w10920w(i) <= estimate_w(i) XOR wire_sincosbitff_w_lg_w_q_range10746w10747w(0);
	END GENERATE loop31;
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7786w8058w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7786w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7868w8141w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7868w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7876w8149w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7876w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7884w8157w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7884w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7892w8165w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7892w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7900w8173w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7900w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7908w8181w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7908w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7916w8189w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7916w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7924w8197w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7924w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7932w8205w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7932w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7940w8213w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7940w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7796w8069w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7796w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7948w8221w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7948w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7956w8229w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7956w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7964w8237w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7964w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7972w8245w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7972w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7980w8253w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7980w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7988w8261w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7988w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7996w8269w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7996w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8004w8277w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8004w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8012w8285w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8012w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8020w8293w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8020w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7804w8077w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7804w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8028w8301w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8028w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8036w8309w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8036w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8044w8317w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8044w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8052w8325w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range8052w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7812w8085w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7812w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7820w8093w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7820w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7828w8101w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7828w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7836w8109w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7836w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7844w8117w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7844w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7852w8125w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7852w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7860w8133w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7860w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8593w8865w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8593w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8675w8948w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8675w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8683w8956w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8683w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8691w8964w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8691w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8699w8972w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8699w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8707w8980w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8707w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8715w8988w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8715w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8723w8996w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8723w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8731w9004w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8731w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8739w9012w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8739w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8747w9020w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8747w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8603w8876w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8603w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8755w9028w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8755w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8763w9036w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8763w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8771w9044w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8771w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8779w9052w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8779w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8787w9060w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8787w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8795w9068w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8795w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8803w9076w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8803w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8811w9084w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8811w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8819w9092w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8819w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8827w9100w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8827w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8611w8884w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8611w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8835w9108w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8835w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8843w9116w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8843w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8851w9124w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8851w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8859w9132w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8859w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8619w8892w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8619w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8627w8900w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8627w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8635w8908w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8635w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8643w8916w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8643w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8651w8924w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8651w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8659w8932w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8659w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8667w8940w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8667w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9395w9667w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9395w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9477w9750w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9477w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9485w9758w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9485w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9493w9766w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9493w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9501w9774w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9501w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9509w9782w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9509w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9517w9790w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9517w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9525w9798w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9525w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9533w9806w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9533w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9541w9814w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9541w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9549w9822w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9549w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9405w9678w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9405w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9557w9830w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9557w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9565w9838w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9565w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9573w9846w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9573w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9581w9854w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9581w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9589w9862w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9589w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9597w9870w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9597w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9605w9878w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9605w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9613w9886w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9613w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9621w9894w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9621w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9629w9902w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9629w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9413w9686w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9413w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9637w9910w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9637w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9645w9918w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9645w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9653w9926w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9653w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9661w9934w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9661w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9421w9694w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9421w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9429w9702w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9429w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9437w9710w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9437w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9445w9718w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9445w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9453w9726w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9453w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9461w9734w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9461w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9469w9742w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range9469w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10192w10464w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10192w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10274w10547w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10274w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10282w10555w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10282w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10290w10563w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10290w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10298w10571w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10298w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10306w10579w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10306w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10314w10587w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10314w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10322w10595w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10322w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10330w10603w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10330w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10338w10611w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10338w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10346w10619w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10346w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10202w10475w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10202w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10354w10627w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10354w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10362w10635w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10362w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10370w10643w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10370w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10378w10651w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10378w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10386w10659w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10386w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10394w10667w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10394w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10402w10675w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10402w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10410w10683w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10410w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10418w10691w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10418w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10426w10699w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10426w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10210w10483w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10210w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10434w10707w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10434w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10442w10715w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10442w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10450w10723w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10450w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10458w10731w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10458w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10218w10491w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10218w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10226w10499w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10226w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10234w10507w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10234w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10242w10515w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10242w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10250w10523w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10250w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10258w10531w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10258w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10266w10539w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range10266w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1150w1422w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1150w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1232w1505w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1232w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1240w1513w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1240w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1248w1521w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1248w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1256w1529w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1256w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1264w1537w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1264w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1272w1545w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1272w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1280w1553w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1280w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1288w1561w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1288w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1296w1569w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1296w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1304w1577w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1304w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1160w1433w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1160w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1312w1585w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1312w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1320w1593w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1320w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1328w1601w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1328w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1336w1609w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1336w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1344w1617w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1344w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1352w1625w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1352w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1360w1633w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1360w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1368w1641w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1368w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1376w1649w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1376w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1384w1657w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1384w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1168w1441w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1168w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1392w1665w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1392w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1400w1673w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1400w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1408w1681w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1408w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1416w1689w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1416w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1176w1449w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1176w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1184w1457w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1184w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1192w1465w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1192w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1200w1473w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1200w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1208w1481w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1208w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1216w1489w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1216w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1224w1497w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1224w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1997w2269w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1997w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2079w2352w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2079w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2087w2360w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2087w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2095w2368w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2095w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2103w2376w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2103w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2111w2384w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2111w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2119w2392w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2119w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2127w2400w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2127w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2135w2408w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2135w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2143w2416w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2143w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2151w2424w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2151w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2007w2280w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2007w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2159w2432w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2159w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2167w2440w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2167w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2175w2448w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2175w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2183w2456w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2183w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2191w2464w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2191w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2199w2472w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2199w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2207w2480w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2207w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2215w2488w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2215w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2223w2496w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2223w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2231w2504w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2231w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2015w2288w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2015w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2239w2512w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2239w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2247w2520w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2247w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2255w2528w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2255w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2263w2536w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2263w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2023w2296w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2023w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2031w2304w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2031w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2039w2312w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2039w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2047w2320w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2047w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2055w2328w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2055w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2063w2336w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2063w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2071w2344w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2071w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2839w3111w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2839w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2921w3194w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2921w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2929w3202w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2929w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2937w3210w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2937w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2945w3218w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2945w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2953w3226w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2953w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2961w3234w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2961w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2969w3242w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2969w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2977w3250w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2977w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2985w3258w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2985w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2993w3266w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2993w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2849w3122w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2849w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3001w3274w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3001w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3009w3282w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3009w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3017w3290w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3017w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3025w3298w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3025w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3033w3306w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3033w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3041w3314w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3041w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3049w3322w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3049w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3057w3330w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3057w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3065w3338w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3065w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3073w3346w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3073w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2857w3130w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2857w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3081w3354w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3081w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3089w3362w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3089w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3097w3370w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3097w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3105w3378w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range3105w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2865w3138w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2865w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2873w3146w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2873w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2881w3154w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2881w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2889w3162w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2889w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2897w3170w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2897w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2905w3178w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2905w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2913w3186w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2913w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3676w3948w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3676w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3758w4031w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3758w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3766w4039w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3766w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3774w4047w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3774w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3782w4055w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3782w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3790w4063w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3790w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3798w4071w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3798w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3806w4079w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3806w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3814w4087w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3814w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3822w4095w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3822w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3830w4103w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3830w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3686w3959w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3686w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3838w4111w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3838w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3846w4119w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3846w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3854w4127w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3854w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3862w4135w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3862w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3870w4143w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3870w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3878w4151w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3878w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3886w4159w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3886w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3894w4167w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3894w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3902w4175w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3902w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3910w4183w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3910w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3694w3967w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3694w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3918w4191w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3918w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3926w4199w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3926w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3934w4207w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3934w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3942w4215w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3942w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3702w3975w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3702w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3710w3983w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3710w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3718w3991w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3718w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3726w3999w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3726w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3734w4007w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3734w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3742w4015w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3742w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3750w4023w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3750w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4508w4780w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4508w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4590w4863w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4590w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4598w4871w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4598w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4606w4879w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4606w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4614w4887w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4614w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4622w4895w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4622w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4630w4903w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4630w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4638w4911w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4638w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4646w4919w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4646w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4654w4927w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4654w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4662w4935w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4662w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4518w4791w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4518w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4670w4943w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4670w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4678w4951w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4678w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4686w4959w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4686w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4694w4967w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4694w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4702w4975w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4702w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4710w4983w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4710w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4718w4991w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4718w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4726w4999w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4726w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4734w5007w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4734w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4742w5015w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4742w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4526w4799w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4526w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4750w5023w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4750w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4758w5031w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4758w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4766w5039w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4766w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4774w5047w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4774w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4534w4807w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4534w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4542w4815w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4542w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4550w4823w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4550w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4558w4831w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4558w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4566w4839w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4566w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4574w4847w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4574w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4582w4855w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4582w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5335w5607w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5335w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5417w5690w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5417w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5425w5698w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5425w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5433w5706w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5433w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5441w5714w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5441w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5449w5722w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5449w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5457w5730w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5457w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5465w5738w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5465w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5473w5746w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5473w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5481w5754w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5481w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5489w5762w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5489w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5345w5618w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5345w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5497w5770w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5497w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5505w5778w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5505w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5513w5786w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5513w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5521w5794w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5521w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5529w5802w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5529w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5537w5810w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5537w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5545w5818w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5545w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5553w5826w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5553w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5561w5834w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5561w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5569w5842w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5569w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5353w5626w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5353w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5577w5850w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5577w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5585w5858w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5585w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5593w5866w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5593w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5601w5874w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5601w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5361w5634w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5361w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5369w5642w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5369w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5377w5650w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5377w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5385w5658w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5385w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5393w5666w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5393w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5401w5674w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5401w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5409w5682w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5409w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6157w6429w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6157w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6239w6512w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6239w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6247w6520w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6247w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6255w6528w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6255w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6263w6536w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6263w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6271w6544w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6271w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6279w6552w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6279w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6287w6560w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6287w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6295w6568w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6295w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6303w6576w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6303w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6311w6584w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6311w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6167w6440w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6167w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6319w6592w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6319w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6327w6600w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6327w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6335w6608w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6335w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6343w6616w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6343w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6351w6624w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6351w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6359w6632w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6359w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6367w6640w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6367w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6375w6648w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6375w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6383w6656w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6383w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6391w6664w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6391w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6175w6448w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6175w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6399w6672w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6399w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6407w6680w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6407w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6415w6688w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6415w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6423w6696w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6423w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6183w6456w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6183w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6191w6464w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6191w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6199w6472w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6199w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6207w6480w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6207w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6215w6488w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6215w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6223w6496w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6223w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6231w6504w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range6231w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6974w7246w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6974w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7056w7329w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7056w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7064w7337w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7064w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7072w7345w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7072w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7080w7353w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7080w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7088w7361w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7088w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7096w7369w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7096w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7104w7377w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7104w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7112w7385w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7112w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7120w7393w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7120w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7128w7401w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7128w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6984w7257w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6984w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7136w7409w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7136w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7144w7417w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7144w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7152w7425w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7152w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7160w7433w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7160w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7168w7441w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7168w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7176w7449w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7176w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7184w7457w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7184w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7192w7465w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7192w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7200w7473w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7200w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7208w7481w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7208w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6992w7265w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6992w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7216w7489w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7216w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7224w7497w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7224w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7232w7505w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7232w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7240w7513w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7240w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7000w7273w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7000w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7008w7281w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7008w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7016w7289w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7016w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7024w7297w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7024w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7032w7305w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7032w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7040w7313w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7040w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7048w7321w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range7048w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7791w8061w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7791w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7872w8143w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7872w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7880w8151w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7880w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7888w8159w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7888w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7896w8167w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7896w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7904w8175w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7904w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7912w8183w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7912w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7920w8191w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7920w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7928w8199w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7928w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7936w8207w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7936w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7944w8215w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7944w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7800w8071w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7800w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7952w8223w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7952w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7960w8231w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7960w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7968w8239w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7968w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7976w8247w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7976w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7984w8255w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7984w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7992w8263w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7992w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8000w8271w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8000w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8008w8279w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8008w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8016w8287w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8016w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8024w8295w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8024w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7808w8079w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7808w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8032w8303w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8032w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8040w8311w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8040w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8048w8319w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8048w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8056w8327w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range8056w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7816w8087w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7816w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7824w8095w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7824w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7832w8103w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7832w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7840w8111w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7840w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7848w8119w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7848w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7856w8127w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7856w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7864w8135w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7864w(0) XOR wire_z_pipeff_9_w_q_range8057w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8598w8868w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8598w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8679w8950w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8679w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8687w8958w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8687w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8695w8966w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8695w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8703w8974w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8703w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8711w8982w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8711w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8719w8990w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8719w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8727w8998w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8727w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8735w9006w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8735w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8743w9014w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8743w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8751w9022w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8751w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8607w8878w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8607w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8759w9030w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8759w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8767w9038w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8767w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8775w9046w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8775w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8783w9054w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8783w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8791w9062w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8791w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8799w9070w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8799w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8807w9078w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8807w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8815w9086w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8815w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8823w9094w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8823w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8831w9102w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8831w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8615w8886w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8615w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8839w9110w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8839w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8847w9118w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8847w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8855w9126w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8855w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8863w9134w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8863w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8623w8894w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8623w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8631w8902w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8631w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8639w8910w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8639w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8647w8918w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8647w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8655w8926w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8655w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8663w8934w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8663w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8671w8942w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8671w(0) XOR wire_z_pipeff_10_w_q_range8864w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9400w9670w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9400w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9481w9752w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9481w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9489w9760w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9489w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9497w9768w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9497w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9505w9776w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9505w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9513w9784w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9513w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9521w9792w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9521w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9529w9800w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9529w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9537w9808w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9537w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9545w9816w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9545w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9553w9824w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9553w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9409w9680w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9409w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9561w9832w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9561w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9569w9840w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9569w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9577w9848w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9577w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9585w9856w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9585w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9593w9864w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9593w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9601w9872w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9601w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9609w9880w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9609w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9617w9888w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9617w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9625w9896w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9625w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9633w9904w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9633w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9417w9688w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9417w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9641w9912w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9641w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9649w9920w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9649w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9657w9928w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9657w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9665w9936w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9665w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9425w9696w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9425w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9433w9704w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9433w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9441w9712w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9441w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9449w9720w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9449w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9457w9728w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9457w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9465w9736w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9465w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9473w9744w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range9473w(0) XOR wire_z_pipeff_11_w_q_range9666w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10197w10467w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10197w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10278w10549w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10278w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10286w10557w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10286w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10294w10565w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10294w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10302w10573w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10302w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10310w10581w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10310w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10318w10589w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10318w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10326w10597w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10326w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10334w10605w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10334w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10342w10613w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10342w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10350w10621w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10350w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10206w10477w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10206w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10358w10629w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10358w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10366w10637w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10366w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10374w10645w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10374w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10382w10653w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10382w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10390w10661w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10390w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10398w10669w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10398w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10406w10677w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10406w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10414w10685w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10414w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10422w10693w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10422w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10430w10701w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10430w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10214w10485w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10214w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10438w10709w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10438w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10446w10717w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10446w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10454w10725w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10454w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10462w10733w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10462w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10222w10493w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10222w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10230w10501w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10230w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10238w10509w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10238w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10246w10517w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10246w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10254w10525w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10254w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10262w10533w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10262w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10270w10541w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range10270w(0) XOR wire_z_pipeff_12_w_q_range10463w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1155w1425w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1155w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1236w1507w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1236w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1244w1515w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1244w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1252w1523w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1252w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1260w1531w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1260w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1268w1539w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1268w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1276w1547w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1276w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1284w1555w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1284w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1292w1563w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1292w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1300w1571w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1300w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1308w1579w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1308w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1164w1435w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1164w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1316w1587w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1316w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1324w1595w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1324w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1332w1603w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1332w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1340w1611w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1340w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1348w1619w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1348w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1356w1627w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1356w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1364w1635w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1364w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1372w1643w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1372w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1380w1651w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1380w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1388w1659w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1388w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1172w1443w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1172w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1396w1667w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1396w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1404w1675w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1404w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1412w1683w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1412w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1420w1691w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1420w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1180w1451w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1180w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1188w1459w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1188w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1196w1467w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1196w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1204w1475w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1204w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1212w1483w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1212w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1220w1491w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1220w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1228w1499w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1228w(0) XOR wire_z_pipeff_1_w_q_range1421w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2002w2272w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2002w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2083w2354w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2083w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2091w2362w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2091w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2099w2370w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2099w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2107w2378w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2107w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2115w2386w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2115w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2123w2394w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2123w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2131w2402w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2131w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2139w2410w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2139w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2147w2418w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2147w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2155w2426w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2155w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2011w2282w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2011w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2163w2434w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2163w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2171w2442w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2171w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2179w2450w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2179w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2187w2458w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2187w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2195w2466w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2195w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2203w2474w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2203w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2211w2482w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2211w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2219w2490w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2219w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2227w2498w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2227w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2235w2506w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2235w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2019w2290w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2019w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2243w2514w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2243w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2251w2522w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2251w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2259w2530w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2259w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2267w2538w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2267w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2027w2298w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2027w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2035w2306w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2035w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2043w2314w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2043w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2051w2322w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2051w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2059w2330w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2059w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2067w2338w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2067w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2075w2346w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2075w(0) XOR wire_z_pipeff_2_w_q_range2268w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2844w3114w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2844w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2925w3196w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2925w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2933w3204w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2933w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2941w3212w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2941w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2949w3220w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2949w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2957w3228w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2957w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2965w3236w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2965w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2973w3244w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2973w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2981w3252w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2981w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2989w3260w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2989w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2997w3268w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2997w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2853w3124w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2853w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3005w3276w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3005w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3013w3284w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3013w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3021w3292w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3021w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3029w3300w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3029w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3037w3308w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3037w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3045w3316w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3045w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3053w3324w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3053w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3061w3332w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3061w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3069w3340w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3069w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3077w3348w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3077w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2861w3132w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2861w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3085w3356w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3085w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3093w3364w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3093w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3101w3372w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3101w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3109w3380w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range3109w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2869w3140w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2869w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2877w3148w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2877w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2885w3156w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2885w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2893w3164w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2893w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2901w3172w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2901w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2909w3180w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2909w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2917w3188w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2917w(0) XOR wire_z_pipeff_3_w_q_range3110w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3681w3951w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3681w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3762w4033w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3762w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3770w4041w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3770w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3778w4049w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3778w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3786w4057w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3786w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3794w4065w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3794w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3802w4073w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3802w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3810w4081w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3810w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3818w4089w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3818w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3826w4097w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3826w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3834w4105w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3834w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3690w3961w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3690w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3842w4113w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3842w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3850w4121w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3850w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3858w4129w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3858w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3866w4137w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3866w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3874w4145w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3874w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3882w4153w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3882w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3890w4161w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3890w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3898w4169w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3898w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3906w4177w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3906w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3914w4185w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3914w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3698w3969w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3698w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3922w4193w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3922w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3930w4201w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3930w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3938w4209w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3938w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3946w4217w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3946w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3706w3977w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3706w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3714w3985w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3714w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3722w3993w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3722w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3730w4001w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3730w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3738w4009w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3738w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3746w4017w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3746w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3754w4025w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3754w(0) XOR wire_z_pipeff_4_w_q_range3947w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4513w4783w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4513w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4594w4865w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4594w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4602w4873w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4602w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4610w4881w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4610w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4618w4889w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4618w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4626w4897w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4626w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4634w4905w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4634w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4642w4913w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4642w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4650w4921w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4650w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4658w4929w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4658w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4666w4937w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4666w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4522w4793w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4522w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4674w4945w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4674w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4682w4953w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4682w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4690w4961w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4690w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4698w4969w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4698w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4706w4977w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4706w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4714w4985w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4714w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4722w4993w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4722w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4730w5001w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4730w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4738w5009w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4738w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4746w5017w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4746w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4530w4801w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4530w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4754w5025w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4754w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4762w5033w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4762w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4770w5041w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4770w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4778w5049w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4778w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4538w4809w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4538w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4546w4817w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4546w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4554w4825w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4554w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4562w4833w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4562w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4570w4841w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4570w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4578w4849w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4578w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4586w4857w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4586w(0) XOR wire_z_pipeff_5_w_q_range4779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5340w5610w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5340w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5421w5692w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5421w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5429w5700w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5429w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5437w5708w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5437w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5445w5716w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5445w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5453w5724w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5453w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5461w5732w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5461w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5469w5740w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5469w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5477w5748w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5477w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5485w5756w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5485w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5493w5764w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5493w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5349w5620w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5349w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5501w5772w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5501w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5509w5780w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5509w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5517w5788w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5517w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5525w5796w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5525w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5533w5804w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5533w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5541w5812w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5541w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5549w5820w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5549w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5557w5828w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5557w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5565w5836w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5565w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5573w5844w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5573w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5357w5628w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5357w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5581w5852w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5581w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5589w5860w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5589w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5597w5868w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5597w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5605w5876w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5605w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5365w5636w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5365w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5373w5644w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5373w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5381w5652w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5381w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5389w5660w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5389w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5397w5668w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5397w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5405w5676w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5405w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5413w5684w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5413w(0) XOR wire_z_pipeff_6_w_q_range5606w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6162w6432w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6162w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6243w6514w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6243w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6251w6522w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6251w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6259w6530w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6259w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6267w6538w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6267w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6275w6546w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6275w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6283w6554w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6283w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6291w6562w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6291w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6299w6570w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6299w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6307w6578w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6307w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6315w6586w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6315w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6171w6442w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6171w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6323w6594w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6323w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6331w6602w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6331w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6339w6610w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6339w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6347w6618w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6347w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6355w6626w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6355w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6363w6634w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6363w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6371w6642w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6371w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6379w6650w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6379w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6387w6658w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6387w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6395w6666w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6395w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6179w6450w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6179w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6403w6674w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6403w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6411w6682w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6411w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6419w6690w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6419w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6427w6698w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6427w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6187w6458w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6187w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6195w6466w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6195w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6203w6474w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6203w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6211w6482w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6211w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6219w6490w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6219w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6227w6498w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6227w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6235w6506w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range6235w(0) XOR wire_z_pipeff_7_w_q_range6428w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6979w7249w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6979w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7060w7331w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7060w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7068w7339w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7068w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7076w7347w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7076w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7084w7355w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7084w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7092w7363w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7092w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7100w7371w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7100w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7108w7379w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7108w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7116w7387w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7116w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7124w7395w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7124w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7132w7403w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7132w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6988w7259w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6988w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7140w7411w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7140w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7148w7419w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7148w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7156w7427w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7156w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7164w7435w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7164w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7172w7443w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7172w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7180w7451w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7180w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7188w7459w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7188w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7196w7467w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7196w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7204w7475w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7204w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7212w7483w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7212w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6996w7267w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6996w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7220w7491w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7220w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7228w7499w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7228w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7236w7507w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7236w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7244w7515w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7244w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7004w7275w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7004w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7012w7283w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7012w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7020w7291w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7020w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7028w7299w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7028w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7036w7307w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7036w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7044w7315w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7044w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7052w7323w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range7052w(0) XOR wire_z_pipeff_8_w_q_range7245w(0);
	atannode_0_w <= wire_cata_0_cordic_atan_arctan;
	atannode_10_w <= wire_cata_10_cordic_atan_arctan;
	atannode_11_w <= wire_cata_11_cordic_atan_arctan;
	atannode_12_w <= wire_cata_12_cordic_atan_arctan;
	atannode_1_w <= wire_cata_1_cordic_atan_arctan;
	atannode_2_w <= wire_cata_2_cordic_atan_arctan;
	atannode_3_w <= wire_cata_3_cordic_atan_arctan;
	atannode_4_w <= wire_cata_4_cordic_atan_arctan;
	atannode_5_w <= wire_cata_5_cordic_atan_arctan;
	atannode_6_w <= wire_cata_6_cordic_atan_arctan;
	atannode_7_w <= wire_cata_7_cordic_atan_arctan;
	atannode_8_w <= wire_cata_8_cordic_atan_arctan;
	atannode_9_w <= wire_cata_9_cordic_atan_arctan;
	delay_input_w <= (wire_x_pipeff_13_w_lg_q10744w OR wire_y_pipeff_13_w_lg_q10743w);
	delay_pipe_w <= cdaff_2;
	estimate_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10909w10917w10918w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10904w10914w10915w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10899w10911w10912w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10894w10906w10907w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10889w10901w10902w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10884w10896w10897w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10879w10891w10892w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10874w10886w10887w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10869w10881w10882w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10864w10876w10877w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10859w10871w10872w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10854w10866w10867w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10849w10861w10862w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10844w10856w10857w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10839w10851w10852w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10834w10846w10847w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10829w10841w10842w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10824w10836w10837w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10819w10831w10832w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10814w10826w10827w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10809w10821w10822w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10804w10816w10817w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10799w10811w10812w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10794w10806w10807w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10789w10801w10802w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10784w10796w10797w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10779w10791w10792w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10774w10786w10787w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10769w10781w10782w
 & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10764w10776w10777w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10758w10771w10772w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10750w10766w10767w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10760w10761w10762w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10753w10754w10755w);
	indexpointnum_w <= (OTHERS => '0');
	multiplier_input_w <= (wire_x_pipeff_13_w_lg_q10741w OR wire_y_pipeff_13_w_lg_q10740w);
	multipliernode_w <= wire_cmx_result;
	post_estimate_w <= wire_ccc_cordic_m_w_lg_estimate_w10920w;
	pre_estimate_w <= multipliernode_w(65 DOWNTO 32);
	radians_load_node_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_radians_range573w576w577w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range568w571w572w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range563w566w567w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range558w561w562w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range553w556w557w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range548w551w552w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range543w546w547w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range538w541w542w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range533w536w537w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range528w531w532w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range523w526w527w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range518w521w522w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range513w516w517w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range508w511w512w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range503w506w507w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range498w501w502w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range493w496w497w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range488w491w492w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range483w486w487w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range478w481w482w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range473w476w477w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range468w471w472w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range463w466w467w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range458w461w462w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range453w456w457w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range448w451w452w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range443w446w447w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range438w441w442w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range433w436w437w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range428w431w432w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range423w426w427w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range418w421w422w & wire_ccc_cordic_m_w_lg_w_radians_range415w417w & wire_ccc_cordic_m_w_lg_w_radians_range410w413w);
	sincos <= sincosff;
	startindex_w <= wire_ccc_cordic_m_w_lg_indexpointnum_w409w;
	x_pipenode_10_w <= wire_x_pipenode_10_add_result;
	x_pipenode_11_w <= wire_x_pipenode_11_add_result;
	x_pipenode_12_w <= wire_x_pipenode_12_add_result;
	x_pipenode_13_w <= wire_x_pipenode_13_add_result;
	x_pipenode_2_w <= wire_x_pipenode_2_add_result;
	x_pipenode_3_w <= wire_x_pipenode_3_add_result;
	x_pipenode_4_w <= wire_x_pipenode_4_add_result;
	x_pipenode_5_w <= wire_x_pipenode_5_add_result;
	x_pipenode_6_w <= wire_x_pipenode_6_add_result;
	x_pipenode_7_w <= wire_x_pipenode_7_add_result;
	x_pipenode_8_w <= wire_x_pipenode_8_add_result;
	x_pipenode_9_w <= wire_x_pipenode_9_add_result;
	x_prenode_10_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7542w8050w8051w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7540w8042w8043w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7538w8034w8035w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7536w8026w8027w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7534w8018w8019w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7532w8010w8011w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7530w8002w8003w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7528w7994w7995w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7523w7986w7987w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7711w7978w7979w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7707w7970w7971w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7701w7962w7963w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7695w7954w7955w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7689w7946w7947w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7683w7938w7939w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7677w7930w7931w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7671w7922w7923w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7665w7914w7915w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7659w7906w7907w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7653w7898w7899w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7647w7890w7891w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7641w7882w7883w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7635w7874w7875w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7629w7866w7867w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7623w7858w7859w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7617w7850w7851w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7611w7842w7843w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7605w7834w7835w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7599w7826w7827w
 & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7593w7818w7819w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7587w7810w7811w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7581w7802w7803w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7575w7794w7795w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7570w7784w7785w);
	x_prenode_11_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8356w8857w8858w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8354w8849w8850w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8352w8841w8842w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8350w8833w8834w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8348w8825w8826w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8346w8817w8818w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8344w8809w8810w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8342w8801w8802w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8340w8793w8794w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8335w8785w8786w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8521w8777w8778w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8517w8769w8770w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8511w8761w8762w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8505w8753w8754w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8499w8745w8746w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8493w8737w8738w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8487w8729w8730w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8481w8721w8722w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8475w8713w8714w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8469w8705w8706w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8463w8697w8698w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8457w8689w8690w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8451w8681w8682w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8445w8673w8674w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8439w8665w8666w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8433w8657w8658w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8427w8649w8650w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8421w8641w8642w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8415w8633w8634w
 & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8409w8625w8626w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8403w8617w8618w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8397w8609w8610w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8391w8601w8602w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range8386w8591w8592w);
	x_prenode_12_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9165w9659w9660w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9163w9651w9652w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9161w9643w9644w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9159w9635w9636w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9157w9627w9628w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9155w9619w9620w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9153w9611w9612w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9151w9603w9604w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9149w9595w9596w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9147w9587w9588w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9142w9579w9580w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9326w9571w9572w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9322w9563w9564w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9316w9555w9556w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9310w9547w9548w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9304w9539w9540w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9298w9531w9532w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9292w9523w9524w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9286w9515w9516w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9280w9507w9508w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9274w9499w9500w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9268w9491w9492w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9262w9483w9484w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9256w9475w9476w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9250w9467w9468w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9244w9459w9460w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9238w9451w9452w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9232w9443w9444w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9226w9435w9436w
 & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9220w9427w9428w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9214w9419w9420w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9208w9411w9412w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9202w9403w9404w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range9197w9393w9394w);
	x_prenode_13_w <= ( wire_ccc_cordic_m_w10457w & wire_ccc_cordic_m_w10449w & wire_ccc_cordic_m_w10441w & wire_ccc_cordic_m_w10433w & wire_ccc_cordic_m_w10425w & wire_ccc_cordic_m_w10417w & wire_ccc_cordic_m_w10409w & wire_ccc_cordic_m_w10401w & wire_ccc_cordic_m_w10393w & wire_ccc_cordic_m_w10385w & wire_ccc_cordic_m_w10377w & wire_ccc_cordic_m_w10369w & wire_ccc_cordic_m_w10361w & wire_ccc_cordic_m_w10353w & wire_ccc_cordic_m_w10345w & wire_ccc_cordic_m_w10337w & wire_ccc_cordic_m_w10329w & wire_ccc_cordic_m_w10321w & wire_ccc_cordic_m_w10313w & wire_ccc_cordic_m_w10305w & wire_ccc_cordic_m_w10297w & wire_ccc_cordic_m_w10289w & wire_ccc_cordic_m_w10281w & wire_ccc_cordic_m_w10273w & wire_ccc_cordic_m_w10265w & wire_ccc_cordic_m_w10257w & wire_ccc_cordic_m_w10249w & wire_ccc_cordic_m_w10241w & wire_ccc_cordic_m_w10233w & wire_ccc_cordic_m_w10225w & wire_ccc_cordic_m_w10217w & wire_ccc_cordic_m_w10209w & wire_ccc_cordic_m_w10201w & wire_ccc_cordic_m_w10191w);
	x_prenode_2_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range847w1414w1415w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1051w1406w1407w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1047w1398w1399w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1041w1390w1391w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1035w1382w1383w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1029w1374w1375w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1023w1366w1367w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1017w1358w1359w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1011w1350w1351w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range1005w1342w1343w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range999w1334w1335w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range993w1326w1327w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range987w1318w1319w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range981w1310w1311w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range975w1302w1303w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range969w1294w1295w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range963w1286w1287w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range957w1278w1279w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range951w1270w1271w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range945w1262w1263w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range939w1254w1255w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range933w1246w1247w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range927w1238w1239w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range921w1230w1231w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range915w1222w1223w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range909w1214w1215w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range903w1206w1207w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range897w1198w1199w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range891w1190w1191w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range885w1182w1183w
 & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range879w1174w1175w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range873w1166w1167w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range867w1158w1159w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range862w1148w1149w);
	x_prenode_3_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1704w2261w2262w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1699w2253w2254w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1901w2245w2246w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1897w2237w2238w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1891w2229w2230w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1885w2221w2222w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1879w2213w2214w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1873w2205w2206w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1867w2197w2198w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1861w2189w2190w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1855w2181w2182w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1849w2173w2174w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1843w2165w2166w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1837w2157w2158w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1831w2149w2150w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1825w2141w2142w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1819w2133w2134w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1813w2125w2126w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1807w2117w2118w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1801w2109w2110w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1795w2101w2102w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1789w2093w2094w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1783w2085w2086w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1777w2077w2078w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1771w2069w2070w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1765w2061w2062w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1759w2053w2054w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1753w2045w2046w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1747w2037w2038w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1741w2029w2030w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1735w2021w2022w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1729w2013w2014w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1723w2005w2006w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1718w1995w1996w);
	x_prenode_4_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2553w3103w3104w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2551w3095w3096w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2546w3087w3088w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2746w3079w3080w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2742w3071w3072w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2736w3063w3064w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2730w3055w3056w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2724w3047w3048w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2718w3039w3040w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2712w3031w3032w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2706w3023w3024w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2700w3015w3016w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2694w3007w3008w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2688w2999w3000w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2682w2991w2992w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2676w2983w2984w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2670w2975w2976w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2664w2967w2968w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2658w2959w2960w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2652w2951w2952w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2646w2943w2944w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2640w2935w2936w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2634w2927w2928w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2628w2919w2920w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2622w2911w2912w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2616w2903w2904w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2610w2895w2896w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2604w2887w2888w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2598w2879w2880w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2592w2871w2872w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2586w2863w2864w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2580w2855w2856w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2574w2847w2848w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2569w2837w2838w);
	x_prenode_5_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3397w3940w3941w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3395w3932w3933w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3393w3924w3925w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3388w3916w3917w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3586w3908w3909w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3582w3900w3901w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3576w3892w3893w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3570w3884w3885w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3564w3876w3877w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3558w3868w3869w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3552w3860w3861w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3546w3852w3853w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3540w3844w3845w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3534w3836w3837w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3528w3828w3829w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3522w3820w3821w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3516w3812w3813w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3510w3804w3805w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3504w3796w3797w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3498w3788w3789w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3492w3780w3781w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3486w3772w3773w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3480w3764w3765w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3474w3756w3757w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3468w3748w3749w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3462w3740w3741w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3456w3732w3733w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3450w3724w3725w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3444w3716w3717w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3438w3708w3709w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3432w3700w3701w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3426w3692w3693w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3420w3684w3685w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3415w3674w3675w);
	x_prenode_6_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4236w4772w4773w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4234w4764w4765w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4232w4756w4757w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4230w4748w4749w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4225w4740w4741w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4421w4732w4733w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4417w4724w4725w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4411w4716w4717w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4405w4708w4709w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4399w4700w4701w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4393w4692w4693w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4387w4684w4685w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4381w4676w4677w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4375w4668w4669w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4369w4660w4661w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4363w4652w4653w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4357w4644w4645w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4351w4636w4637w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4345w4628w4629w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4339w4620w4621w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4333w4612w4613w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4327w4604w4605w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4321w4596w4597w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4315w4588w4589w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4309w4580w4581w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4303w4572w4573w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4297w4564w4565w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4291w4556w4557w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4285w4548w4549w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4279w4540w4541w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4273w4532w4533w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4267w4524w4525w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4261w4516w4517w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4256w4506w4507w);
	x_prenode_7_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5070w5599w5600w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5068w5591w5592w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5066w5583w5584w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5064w5575w5576w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5062w5567w5568w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5057w5559w5560w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5251w5551w5552w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5247w5543w5544w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5241w5535w5536w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5235w5527w5528w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5229w5519w5520w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5223w5511w5512w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5217w5503w5504w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5211w5495w5496w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5205w5487w5488w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5199w5479w5480w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5193w5471w5472w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5187w5463w5464w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5181w5455w5456w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5175w5447w5448w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5169w5439w5440w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5163w5431w5432w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5157w5423w5424w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5151w5415w5416w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5145w5407w5408w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5139w5399w5400w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5133w5391w5392w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5127w5383w5384w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5121w5375w5376w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5115w5367w5368w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5109w5359w5360w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5103w5351w5352w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5097w5343w5344w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range5092w5333w5334w);
	x_prenode_8_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5899w6421w6422w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5897w6413w6414w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5895w6405w6406w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5893w6397w6398w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5891w6389w6390w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5889w6381w6382w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5884w6373w6374w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6076w6365w6366w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6072w6357w6358w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6066w6349w6350w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6060w6341w6342w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6054w6333w6334w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6048w6325w6326w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6042w6317w6318w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6036w6309w6310w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6030w6301w6302w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6024w6293w6294w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6018w6285w6286w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6012w6277w6278w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6006w6269w6270w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range6000w6261w6262w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5994w6253w6254w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5988w6245w6246w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5982w6237w6238w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5976w6229w6230w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5970w6221w6222w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5964w6213w6214w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5958w6205w6206w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5952w6197w6198w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5946w6189w6190w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5940w6181w6182w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5934w6173w6174w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5928w6165w6166w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5923w6155w6156w);
	x_prenode_9_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6723w7238w7239w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6721w7230w7231w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6719w7222w7223w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6717w7214w7215w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6715w7206w7207w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6713w7198w7199w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6711w7190w7191w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6706w7182w7183w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6896w7174w7175w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6892w7166w7167w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6886w7158w7159w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6880w7150w7151w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6874w7142w7143w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6868w7134w7135w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6862w7126w7127w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6856w7118w7119w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6850w7110w7111w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6844w7102w7103w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6838w7094w7095w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6832w7086w7087w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6826w7078w7079w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6820w7070w7071w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6814w7062w7063w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6808w7054w7055w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6802w7046w7047w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6796w7038w7039w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6790w7030w7031w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6784w7022w7023w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6778w7014w7015w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6772w7006w7007w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6766w6998w6999w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6760w6990w6991w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6754w6982w6983w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6749w6972w6973w);
	x_prenodeone_10_w <= ( wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7705w7706w & wire_y_pipeff_9_w_lg_w_q_range7699w7700w & wire_y_pipeff_9_w_lg_w_q_range7693w7694w & wire_y_pipeff_9_w_lg_w_q_range7687w7688w & wire_y_pipeff_9_w_lg_w_q_range7681w7682w & wire_y_pipeff_9_w_lg_w_q_range7675w7676w & wire_y_pipeff_9_w_lg_w_q_range7669w7670w & wire_y_pipeff_9_w_lg_w_q_range7663w7664w & wire_y_pipeff_9_w_lg_w_q_range7657w7658w & wire_y_pipeff_9_w_lg_w_q_range7651w7652w & wire_y_pipeff_9_w_lg_w_q_range7645w7646w & wire_y_pipeff_9_w_lg_w_q_range7639w7640w & wire_y_pipeff_9_w_lg_w_q_range7633w7634w & wire_y_pipeff_9_w_lg_w_q_range7627w7628w & wire_y_pipeff_9_w_lg_w_q_range7621w7622w & wire_y_pipeff_9_w_lg_w_q_range7615w7616w & wire_y_pipeff_9_w_lg_w_q_range7609w7610w & wire_y_pipeff_9_w_lg_w_q_range7603w7604w & wire_y_pipeff_9_w_lg_w_q_range7597w7598w & wire_y_pipeff_9_w_lg_w_q_range7591w7592w & wire_y_pipeff_9_w_lg_w_q_range7585w7586w & wire_y_pipeff_9_w_lg_w_q_range7579w7580w & wire_y_pipeff_9_w_lg_w_q_range7573w7574w & wire_y_pipeff_9_w_lg_w_q_range7568w7569w);
	x_prenodeone_11_w <= ( wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8515w8516w & wire_y_pipeff_10_w_lg_w_q_range8509w8510w & wire_y_pipeff_10_w_lg_w_q_range8503w8504w & wire_y_pipeff_10_w_lg_w_q_range8497w8498w & wire_y_pipeff_10_w_lg_w_q_range8491w8492w & wire_y_pipeff_10_w_lg_w_q_range8485w8486w & wire_y_pipeff_10_w_lg_w_q_range8479w8480w & wire_y_pipeff_10_w_lg_w_q_range8473w8474w & wire_y_pipeff_10_w_lg_w_q_range8467w8468w & wire_y_pipeff_10_w_lg_w_q_range8461w8462w & wire_y_pipeff_10_w_lg_w_q_range8455w8456w & wire_y_pipeff_10_w_lg_w_q_range8449w8450w & wire_y_pipeff_10_w_lg_w_q_range8443w8444w & wire_y_pipeff_10_w_lg_w_q_range8437w8438w & wire_y_pipeff_10_w_lg_w_q_range8431w8432w & wire_y_pipeff_10_w_lg_w_q_range8425w8426w & wire_y_pipeff_10_w_lg_w_q_range8419w8420w & wire_y_pipeff_10_w_lg_w_q_range8413w8414w & wire_y_pipeff_10_w_lg_w_q_range8407w8408w & wire_y_pipeff_10_w_lg_w_q_range8401w8402w & wire_y_pipeff_10_w_lg_w_q_range8395w8396w & wire_y_pipeff_10_w_lg_w_q_range8389w8390w & wire_y_pipeff_10_w_lg_w_q_range8384w8385w);
	x_prenodeone_12_w <= ( wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9320w9321w & wire_y_pipeff_11_w_lg_w_q_range9314w9315w & wire_y_pipeff_11_w_lg_w_q_range9308w9309w & wire_y_pipeff_11_w_lg_w_q_range9302w9303w & wire_y_pipeff_11_w_lg_w_q_range9296w9297w & wire_y_pipeff_11_w_lg_w_q_range9290w9291w & wire_y_pipeff_11_w_lg_w_q_range9284w9285w & wire_y_pipeff_11_w_lg_w_q_range9278w9279w & wire_y_pipeff_11_w_lg_w_q_range9272w9273w & wire_y_pipeff_11_w_lg_w_q_range9266w9267w & wire_y_pipeff_11_w_lg_w_q_range9260w9261w & wire_y_pipeff_11_w_lg_w_q_range9254w9255w & wire_y_pipeff_11_w_lg_w_q_range9248w9249w & wire_y_pipeff_11_w_lg_w_q_range9242w9243w & wire_y_pipeff_11_w_lg_w_q_range9236w9237w & wire_y_pipeff_11_w_lg_w_q_range9230w9231w & wire_y_pipeff_11_w_lg_w_q_range9224w9225w & wire_y_pipeff_11_w_lg_w_q_range9218w9219w & wire_y_pipeff_11_w_lg_w_q_range9212w9213w & wire_y_pipeff_11_w_lg_w_q_range9206w9207w & wire_y_pipeff_11_w_lg_w_q_range9200w9201w & wire_y_pipeff_11_w_lg_w_q_range9195w9196w);
	x_prenodeone_13_w <= ( wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range10120w10121w & wire_y_pipeff_12_w_lg_w_q_range10114w10115w & wire_y_pipeff_12_w_lg_w_q_range10108w10109w & wire_y_pipeff_12_w_lg_w_q_range10102w10103w & wire_y_pipeff_12_w_lg_w_q_range10096w10097w & wire_y_pipeff_12_w_lg_w_q_range10090w10091w & wire_y_pipeff_12_w_lg_w_q_range10084w10085w & wire_y_pipeff_12_w_lg_w_q_range10078w10079w & wire_y_pipeff_12_w_lg_w_q_range10072w10073w & wire_y_pipeff_12_w_lg_w_q_range10066w10067w & wire_y_pipeff_12_w_lg_w_q_range10060w10061w & wire_y_pipeff_12_w_lg_w_q_range10054w10055w & wire_y_pipeff_12_w_lg_w_q_range10048w10049w & wire_y_pipeff_12_w_lg_w_q_range10042w10043w & wire_y_pipeff_12_w_lg_w_q_range10036w10037w & wire_y_pipeff_12_w_lg_w_q_range10030w10031w & wire_y_pipeff_12_w_lg_w_q_range10024w10025w & wire_y_pipeff_12_w_lg_w_q_range10018w10019w & wire_y_pipeff_12_w_lg_w_q_range10012w10013w & wire_y_pipeff_12_w_lg_w_q_range10006w10007w & wire_y_pipeff_12_w_lg_w_q_range10001w10002w);
	x_prenodeone_2_w <= ( wire_y_pipeff_1_w_lg_w_q_range845w846w & wire_y_pipeff_1_w_lg_w_q_range845w846w & wire_y_pipeff_1_w_lg_w_q_range1045w1046w & wire_y_pipeff_1_w_lg_w_q_range1039w1040w & wire_y_pipeff_1_w_lg_w_q_range1033w1034w & wire_y_pipeff_1_w_lg_w_q_range1027w1028w & wire_y_pipeff_1_w_lg_w_q_range1021w1022w & wire_y_pipeff_1_w_lg_w_q_range1015w1016w & wire_y_pipeff_1_w_lg_w_q_range1009w1010w & wire_y_pipeff_1_w_lg_w_q_range1003w1004w & wire_y_pipeff_1_w_lg_w_q_range997w998w & wire_y_pipeff_1_w_lg_w_q_range991w992w & wire_y_pipeff_1_w_lg_w_q_range985w986w & wire_y_pipeff_1_w_lg_w_q_range979w980w & wire_y_pipeff_1_w_lg_w_q_range973w974w & wire_y_pipeff_1_w_lg_w_q_range967w968w & wire_y_pipeff_1_w_lg_w_q_range961w962w & wire_y_pipeff_1_w_lg_w_q_range955w956w & wire_y_pipeff_1_w_lg_w_q_range949w950w & wire_y_pipeff_1_w_lg_w_q_range943w944w & wire_y_pipeff_1_w_lg_w_q_range937w938w & wire_y_pipeff_1_w_lg_w_q_range931w932w & wire_y_pipeff_1_w_lg_w_q_range925w926w & wire_y_pipeff_1_w_lg_w_q_range919w920w & wire_y_pipeff_1_w_lg_w_q_range913w914w & wire_y_pipeff_1_w_lg_w_q_range907w908w & wire_y_pipeff_1_w_lg_w_q_range901w902w & wire_y_pipeff_1_w_lg_w_q_range895w896w & wire_y_pipeff_1_w_lg_w_q_range889w890w & wire_y_pipeff_1_w_lg_w_q_range883w884w & wire_y_pipeff_1_w_lg_w_q_range877w878w & wire_y_pipeff_1_w_lg_w_q_range871w872w & wire_y_pipeff_1_w_lg_w_q_range865w866w & wire_y_pipeff_1_w_lg_w_q_range860w861w);
	x_prenodeone_3_w <= ( wire_y_pipeff_2_w_lg_w_q_range1697w1698w & wire_y_pipeff_2_w_lg_w_q_range1697w1698w & wire_y_pipeff_2_w_lg_w_q_range1697w1698w & wire_y_pipeff_2_w_lg_w_q_range1895w1896w & wire_y_pipeff_2_w_lg_w_q_range1889w1890w & wire_y_pipeff_2_w_lg_w_q_range1883w1884w & wire_y_pipeff_2_w_lg_w_q_range1877w1878w & wire_y_pipeff_2_w_lg_w_q_range1871w1872w & wire_y_pipeff_2_w_lg_w_q_range1865w1866w & wire_y_pipeff_2_w_lg_w_q_range1859w1860w & wire_y_pipeff_2_w_lg_w_q_range1853w1854w & wire_y_pipeff_2_w_lg_w_q_range1847w1848w & wire_y_pipeff_2_w_lg_w_q_range1841w1842w & wire_y_pipeff_2_w_lg_w_q_range1835w1836w & wire_y_pipeff_2_w_lg_w_q_range1829w1830w & wire_y_pipeff_2_w_lg_w_q_range1823w1824w & wire_y_pipeff_2_w_lg_w_q_range1817w1818w & wire_y_pipeff_2_w_lg_w_q_range1811w1812w & wire_y_pipeff_2_w_lg_w_q_range1805w1806w & wire_y_pipeff_2_w_lg_w_q_range1799w1800w & wire_y_pipeff_2_w_lg_w_q_range1793w1794w & wire_y_pipeff_2_w_lg_w_q_range1787w1788w & wire_y_pipeff_2_w_lg_w_q_range1781w1782w & wire_y_pipeff_2_w_lg_w_q_range1775w1776w & wire_y_pipeff_2_w_lg_w_q_range1769w1770w & wire_y_pipeff_2_w_lg_w_q_range1763w1764w & wire_y_pipeff_2_w_lg_w_q_range1757w1758w & wire_y_pipeff_2_w_lg_w_q_range1751w1752w & wire_y_pipeff_2_w_lg_w_q_range1745w1746w & wire_y_pipeff_2_w_lg_w_q_range1739w1740w & wire_y_pipeff_2_w_lg_w_q_range1733w1734w & wire_y_pipeff_2_w_lg_w_q_range1727w1728w & wire_y_pipeff_2_w_lg_w_q_range1721w1722w & wire_y_pipeff_2_w_lg_w_q_range1716w1717w);
	x_prenodeone_4_w <= ( wire_y_pipeff_3_w_lg_w_q_range2544w2545w & wire_y_pipeff_3_w_lg_w_q_range2544w2545w & wire_y_pipeff_3_w_lg_w_q_range2544w2545w & wire_y_pipeff_3_w_lg_w_q_range2544w2545w & wire_y_pipeff_3_w_lg_w_q_range2740w2741w & wire_y_pipeff_3_w_lg_w_q_range2734w2735w & wire_y_pipeff_3_w_lg_w_q_range2728w2729w & wire_y_pipeff_3_w_lg_w_q_range2722w2723w & wire_y_pipeff_3_w_lg_w_q_range2716w2717w & wire_y_pipeff_3_w_lg_w_q_range2710w2711w & wire_y_pipeff_3_w_lg_w_q_range2704w2705w & wire_y_pipeff_3_w_lg_w_q_range2698w2699w & wire_y_pipeff_3_w_lg_w_q_range2692w2693w & wire_y_pipeff_3_w_lg_w_q_range2686w2687w & wire_y_pipeff_3_w_lg_w_q_range2680w2681w & wire_y_pipeff_3_w_lg_w_q_range2674w2675w & wire_y_pipeff_3_w_lg_w_q_range2668w2669w & wire_y_pipeff_3_w_lg_w_q_range2662w2663w & wire_y_pipeff_3_w_lg_w_q_range2656w2657w & wire_y_pipeff_3_w_lg_w_q_range2650w2651w & wire_y_pipeff_3_w_lg_w_q_range2644w2645w & wire_y_pipeff_3_w_lg_w_q_range2638w2639w & wire_y_pipeff_3_w_lg_w_q_range2632w2633w & wire_y_pipeff_3_w_lg_w_q_range2626w2627w & wire_y_pipeff_3_w_lg_w_q_range2620w2621w & wire_y_pipeff_3_w_lg_w_q_range2614w2615w & wire_y_pipeff_3_w_lg_w_q_range2608w2609w & wire_y_pipeff_3_w_lg_w_q_range2602w2603w & wire_y_pipeff_3_w_lg_w_q_range2596w2597w & wire_y_pipeff_3_w_lg_w_q_range2590w2591w & wire_y_pipeff_3_w_lg_w_q_range2584w2585w & wire_y_pipeff_3_w_lg_w_q_range2578w2579w & wire_y_pipeff_3_w_lg_w_q_range2572w2573w & wire_y_pipeff_3_w_lg_w_q_range2567w2568w);
	x_prenodeone_5_w <= ( wire_y_pipeff_4_w_lg_w_q_range3386w3387w & wire_y_pipeff_4_w_lg_w_q_range3386w3387w & wire_y_pipeff_4_w_lg_w_q_range3386w3387w & wire_y_pipeff_4_w_lg_w_q_range3386w3387w & wire_y_pipeff_4_w_lg_w_q_range3386w3387w & wire_y_pipeff_4_w_lg_w_q_range3580w3581w & wire_y_pipeff_4_w_lg_w_q_range3574w3575w & wire_y_pipeff_4_w_lg_w_q_range3568w3569w & wire_y_pipeff_4_w_lg_w_q_range3562w3563w & wire_y_pipeff_4_w_lg_w_q_range3556w3557w & wire_y_pipeff_4_w_lg_w_q_range3550w3551w & wire_y_pipeff_4_w_lg_w_q_range3544w3545w & wire_y_pipeff_4_w_lg_w_q_range3538w3539w & wire_y_pipeff_4_w_lg_w_q_range3532w3533w & wire_y_pipeff_4_w_lg_w_q_range3526w3527w & wire_y_pipeff_4_w_lg_w_q_range3520w3521w & wire_y_pipeff_4_w_lg_w_q_range3514w3515w & wire_y_pipeff_4_w_lg_w_q_range3508w3509w & wire_y_pipeff_4_w_lg_w_q_range3502w3503w & wire_y_pipeff_4_w_lg_w_q_range3496w3497w & wire_y_pipeff_4_w_lg_w_q_range3490w3491w & wire_y_pipeff_4_w_lg_w_q_range3484w3485w & wire_y_pipeff_4_w_lg_w_q_range3478w3479w & wire_y_pipeff_4_w_lg_w_q_range3472w3473w & wire_y_pipeff_4_w_lg_w_q_range3466w3467w & wire_y_pipeff_4_w_lg_w_q_range3460w3461w & wire_y_pipeff_4_w_lg_w_q_range3454w3455w & wire_y_pipeff_4_w_lg_w_q_range3448w3449w & wire_y_pipeff_4_w_lg_w_q_range3442w3443w & wire_y_pipeff_4_w_lg_w_q_range3436w3437w & wire_y_pipeff_4_w_lg_w_q_range3430w3431w & wire_y_pipeff_4_w_lg_w_q_range3424w3425w & wire_y_pipeff_4_w_lg_w_q_range3418w3419w & wire_y_pipeff_4_w_lg_w_q_range3413w3414w);
	x_prenodeone_6_w <= ( wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4415w4416w & wire_y_pipeff_5_w_lg_w_q_range4409w4410w & wire_y_pipeff_5_w_lg_w_q_range4403w4404w & wire_y_pipeff_5_w_lg_w_q_range4397w4398w & wire_y_pipeff_5_w_lg_w_q_range4391w4392w & wire_y_pipeff_5_w_lg_w_q_range4385w4386w & wire_y_pipeff_5_w_lg_w_q_range4379w4380w & wire_y_pipeff_5_w_lg_w_q_range4373w4374w & wire_y_pipeff_5_w_lg_w_q_range4367w4368w & wire_y_pipeff_5_w_lg_w_q_range4361w4362w & wire_y_pipeff_5_w_lg_w_q_range4355w4356w & wire_y_pipeff_5_w_lg_w_q_range4349w4350w & wire_y_pipeff_5_w_lg_w_q_range4343w4344w & wire_y_pipeff_5_w_lg_w_q_range4337w4338w & wire_y_pipeff_5_w_lg_w_q_range4331w4332w & wire_y_pipeff_5_w_lg_w_q_range4325w4326w & wire_y_pipeff_5_w_lg_w_q_range4319w4320w & wire_y_pipeff_5_w_lg_w_q_range4313w4314w & wire_y_pipeff_5_w_lg_w_q_range4307w4308w & wire_y_pipeff_5_w_lg_w_q_range4301w4302w & wire_y_pipeff_5_w_lg_w_q_range4295w4296w & wire_y_pipeff_5_w_lg_w_q_range4289w4290w & wire_y_pipeff_5_w_lg_w_q_range4283w4284w & wire_y_pipeff_5_w_lg_w_q_range4277w4278w & wire_y_pipeff_5_w_lg_w_q_range4271w4272w & wire_y_pipeff_5_w_lg_w_q_range4265w4266w & wire_y_pipeff_5_w_lg_w_q_range4259w4260w & wire_y_pipeff_5_w_lg_w_q_range4254w4255w);
	x_prenodeone_7_w <= ( wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5245w5246w & wire_y_pipeff_6_w_lg_w_q_range5239w5240w & wire_y_pipeff_6_w_lg_w_q_range5233w5234w & wire_y_pipeff_6_w_lg_w_q_range5227w5228w & wire_y_pipeff_6_w_lg_w_q_range5221w5222w & wire_y_pipeff_6_w_lg_w_q_range5215w5216w & wire_y_pipeff_6_w_lg_w_q_range5209w5210w & wire_y_pipeff_6_w_lg_w_q_range5203w5204w & wire_y_pipeff_6_w_lg_w_q_range5197w5198w & wire_y_pipeff_6_w_lg_w_q_range5191w5192w & wire_y_pipeff_6_w_lg_w_q_range5185w5186w & wire_y_pipeff_6_w_lg_w_q_range5179w5180w & wire_y_pipeff_6_w_lg_w_q_range5173w5174w & wire_y_pipeff_6_w_lg_w_q_range5167w5168w & wire_y_pipeff_6_w_lg_w_q_range5161w5162w & wire_y_pipeff_6_w_lg_w_q_range5155w5156w & wire_y_pipeff_6_w_lg_w_q_range5149w5150w & wire_y_pipeff_6_w_lg_w_q_range5143w5144w & wire_y_pipeff_6_w_lg_w_q_range5137w5138w & wire_y_pipeff_6_w_lg_w_q_range5131w5132w & wire_y_pipeff_6_w_lg_w_q_range5125w5126w & wire_y_pipeff_6_w_lg_w_q_range5119w5120w & wire_y_pipeff_6_w_lg_w_q_range5113w5114w & wire_y_pipeff_6_w_lg_w_q_range5107w5108w & wire_y_pipeff_6_w_lg_w_q_range5101w5102w & wire_y_pipeff_6_w_lg_w_q_range5095w5096w & wire_y_pipeff_6_w_lg_w_q_range5090w5091w);
	x_prenodeone_8_w <= ( wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range6070w6071w & wire_y_pipeff_7_w_lg_w_q_range6064w6065w & wire_y_pipeff_7_w_lg_w_q_range6058w6059w & wire_y_pipeff_7_w_lg_w_q_range6052w6053w & wire_y_pipeff_7_w_lg_w_q_range6046w6047w & wire_y_pipeff_7_w_lg_w_q_range6040w6041w & wire_y_pipeff_7_w_lg_w_q_range6034w6035w & wire_y_pipeff_7_w_lg_w_q_range6028w6029w & wire_y_pipeff_7_w_lg_w_q_range6022w6023w & wire_y_pipeff_7_w_lg_w_q_range6016w6017w & wire_y_pipeff_7_w_lg_w_q_range6010w6011w & wire_y_pipeff_7_w_lg_w_q_range6004w6005w & wire_y_pipeff_7_w_lg_w_q_range5998w5999w & wire_y_pipeff_7_w_lg_w_q_range5992w5993w & wire_y_pipeff_7_w_lg_w_q_range5986w5987w & wire_y_pipeff_7_w_lg_w_q_range5980w5981w & wire_y_pipeff_7_w_lg_w_q_range5974w5975w & wire_y_pipeff_7_w_lg_w_q_range5968w5969w & wire_y_pipeff_7_w_lg_w_q_range5962w5963w & wire_y_pipeff_7_w_lg_w_q_range5956w5957w & wire_y_pipeff_7_w_lg_w_q_range5950w5951w & wire_y_pipeff_7_w_lg_w_q_range5944w5945w & wire_y_pipeff_7_w_lg_w_q_range5938w5939w & wire_y_pipeff_7_w_lg_w_q_range5932w5933w & wire_y_pipeff_7_w_lg_w_q_range5926w5927w & wire_y_pipeff_7_w_lg_w_q_range5921w5922w);
	x_prenodeone_9_w <= ( wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6890w6891w & wire_y_pipeff_8_w_lg_w_q_range6884w6885w & wire_y_pipeff_8_w_lg_w_q_range6878w6879w & wire_y_pipeff_8_w_lg_w_q_range6872w6873w & wire_y_pipeff_8_w_lg_w_q_range6866w6867w & wire_y_pipeff_8_w_lg_w_q_range6860w6861w & wire_y_pipeff_8_w_lg_w_q_range6854w6855w & wire_y_pipeff_8_w_lg_w_q_range6848w6849w & wire_y_pipeff_8_w_lg_w_q_range6842w6843w & wire_y_pipeff_8_w_lg_w_q_range6836w6837w & wire_y_pipeff_8_w_lg_w_q_range6830w6831w & wire_y_pipeff_8_w_lg_w_q_range6824w6825w & wire_y_pipeff_8_w_lg_w_q_range6818w6819w & wire_y_pipeff_8_w_lg_w_q_range6812w6813w & wire_y_pipeff_8_w_lg_w_q_range6806w6807w & wire_y_pipeff_8_w_lg_w_q_range6800w6801w & wire_y_pipeff_8_w_lg_w_q_range6794w6795w & wire_y_pipeff_8_w_lg_w_q_range6788w6789w & wire_y_pipeff_8_w_lg_w_q_range6782w6783w & wire_y_pipeff_8_w_lg_w_q_range6776w6777w & wire_y_pipeff_8_w_lg_w_q_range6770w6771w & wire_y_pipeff_8_w_lg_w_q_range6764w6765w & wire_y_pipeff_8_w_lg_w_q_range6758w6759w & wire_y_pipeff_8_w_lg_w_q_range6752w6753w & wire_y_pipeff_8_w_lg_w_q_range6747w6748w);
	x_prenodetwo_10_w <= ( wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7521w7522w & wire_y_pipeff_9_w_lg_w_q_range7705w7706w & wire_y_pipeff_9_w_lg_w_q_range7699w7700w & wire_y_pipeff_9_w_lg_w_q_range7693w7694w & wire_y_pipeff_9_w_lg_w_q_range7687w7688w & wire_y_pipeff_9_w_lg_w_q_range7681w7682w & wire_y_pipeff_9_w_lg_w_q_range7675w7676w & wire_y_pipeff_9_w_lg_w_q_range7669w7670w & wire_y_pipeff_9_w_lg_w_q_range7663w7664w & wire_y_pipeff_9_w_lg_w_q_range7657w7658w & wire_y_pipeff_9_w_lg_w_q_range7651w7652w & wire_y_pipeff_9_w_lg_w_q_range7645w7646w & wire_y_pipeff_9_w_lg_w_q_range7639w7640w & wire_y_pipeff_9_w_lg_w_q_range7633w7634w & wire_y_pipeff_9_w_lg_w_q_range7627w7628w & wire_y_pipeff_9_w_lg_w_q_range7621w7622w & wire_y_pipeff_9_w_lg_w_q_range7615w7616w & wire_y_pipeff_9_w_lg_w_q_range7609w7610w & wire_y_pipeff_9_w_lg_w_q_range7603w7604w & wire_y_pipeff_9_w_lg_w_q_range7597w7598w & wire_y_pipeff_9_w_lg_w_q_range7591w7592w & wire_y_pipeff_9_w_lg_w_q_range7585w7586w & wire_y_pipeff_9_w_lg_w_q_range7579w7580w);
	x_prenodetwo_11_w <= ( wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8333w8334w & wire_y_pipeff_10_w_lg_w_q_range8515w8516w & wire_y_pipeff_10_w_lg_w_q_range8509w8510w & wire_y_pipeff_10_w_lg_w_q_range8503w8504w & wire_y_pipeff_10_w_lg_w_q_range8497w8498w & wire_y_pipeff_10_w_lg_w_q_range8491w8492w & wire_y_pipeff_10_w_lg_w_q_range8485w8486w & wire_y_pipeff_10_w_lg_w_q_range8479w8480w & wire_y_pipeff_10_w_lg_w_q_range8473w8474w & wire_y_pipeff_10_w_lg_w_q_range8467w8468w & wire_y_pipeff_10_w_lg_w_q_range8461w8462w & wire_y_pipeff_10_w_lg_w_q_range8455w8456w & wire_y_pipeff_10_w_lg_w_q_range8449w8450w & wire_y_pipeff_10_w_lg_w_q_range8443w8444w & wire_y_pipeff_10_w_lg_w_q_range8437w8438w & wire_y_pipeff_10_w_lg_w_q_range8431w8432w & wire_y_pipeff_10_w_lg_w_q_range8425w8426w & wire_y_pipeff_10_w_lg_w_q_range8419w8420w & wire_y_pipeff_10_w_lg_w_q_range8413w8414w & wire_y_pipeff_10_w_lg_w_q_range8407w8408w & wire_y_pipeff_10_w_lg_w_q_range8401w8402w & wire_y_pipeff_10_w_lg_w_q_range8395w8396w);
	x_prenodetwo_12_w <= ( wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9140w9141w & wire_y_pipeff_11_w_lg_w_q_range9320w9321w & wire_y_pipeff_11_w_lg_w_q_range9314w9315w & wire_y_pipeff_11_w_lg_w_q_range9308w9309w & wire_y_pipeff_11_w_lg_w_q_range9302w9303w & wire_y_pipeff_11_w_lg_w_q_range9296w9297w & wire_y_pipeff_11_w_lg_w_q_range9290w9291w & wire_y_pipeff_11_w_lg_w_q_range9284w9285w & wire_y_pipeff_11_w_lg_w_q_range9278w9279w & wire_y_pipeff_11_w_lg_w_q_range9272w9273w & wire_y_pipeff_11_w_lg_w_q_range9266w9267w & wire_y_pipeff_11_w_lg_w_q_range9260w9261w & wire_y_pipeff_11_w_lg_w_q_range9254w9255w & wire_y_pipeff_11_w_lg_w_q_range9248w9249w & wire_y_pipeff_11_w_lg_w_q_range9242w9243w & wire_y_pipeff_11_w_lg_w_q_range9236w9237w & wire_y_pipeff_11_w_lg_w_q_range9230w9231w & wire_y_pipeff_11_w_lg_w_q_range9224w9225w & wire_y_pipeff_11_w_lg_w_q_range9218w9219w & wire_y_pipeff_11_w_lg_w_q_range9212w9213w & wire_y_pipeff_11_w_lg_w_q_range9206w9207w);
	x_prenodetwo_13_w <= ( wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range9942w9943w & wire_y_pipeff_12_w_lg_w_q_range10120w10121w & wire_y_pipeff_12_w_lg_w_q_range10114w10115w & wire_y_pipeff_12_w_lg_w_q_range10108w10109w & wire_y_pipeff_12_w_lg_w_q_range10102w10103w & wire_y_pipeff_12_w_lg_w_q_range10096w10097w & wire_y_pipeff_12_w_lg_w_q_range10090w10091w & wire_y_pipeff_12_w_lg_w_q_range10084w10085w & wire_y_pipeff_12_w_lg_w_q_range10078w10079w & wire_y_pipeff_12_w_lg_w_q_range10072w10073w & wire_y_pipeff_12_w_lg_w_q_range10066w10067w & wire_y_pipeff_12_w_lg_w_q_range10060w10061w & wire_y_pipeff_12_w_lg_w_q_range10054w10055w & wire_y_pipeff_12_w_lg_w_q_range10048w10049w & wire_y_pipeff_12_w_lg_w_q_range10042w10043w & wire_y_pipeff_12_w_lg_w_q_range10036w10037w & wire_y_pipeff_12_w_lg_w_q_range10030w10031w & wire_y_pipeff_12_w_lg_w_q_range10024w10025w & wire_y_pipeff_12_w_lg_w_q_range10018w10019w & wire_y_pipeff_12_w_lg_w_q_range10012w10013w);
	x_prenodetwo_2_w <= ( wire_y_pipeff_1_w_lg_w_q_range845w846w & wire_y_pipeff_1_w_lg_w_q_range845w846w & wire_y_pipeff_1_w_lg_w_q_range845w846w & wire_y_pipeff_1_w_lg_w_q_range845w846w & wire_y_pipeff_1_w_lg_w_q_range1045w1046w & wire_y_pipeff_1_w_lg_w_q_range1039w1040w & wire_y_pipeff_1_w_lg_w_q_range1033w1034w & wire_y_pipeff_1_w_lg_w_q_range1027w1028w & wire_y_pipeff_1_w_lg_w_q_range1021w1022w & wire_y_pipeff_1_w_lg_w_q_range1015w1016w & wire_y_pipeff_1_w_lg_w_q_range1009w1010w & wire_y_pipeff_1_w_lg_w_q_range1003w1004w & wire_y_pipeff_1_w_lg_w_q_range997w998w & wire_y_pipeff_1_w_lg_w_q_range991w992w & wire_y_pipeff_1_w_lg_w_q_range985w986w & wire_y_pipeff_1_w_lg_w_q_range979w980w & wire_y_pipeff_1_w_lg_w_q_range973w974w & wire_y_pipeff_1_w_lg_w_q_range967w968w & wire_y_pipeff_1_w_lg_w_q_range961w962w & wire_y_pipeff_1_w_lg_w_q_range955w956w & wire_y_pipeff_1_w_lg_w_q_range949w950w & wire_y_pipeff_1_w_lg_w_q_range943w944w & wire_y_pipeff_1_w_lg_w_q_range937w938w & wire_y_pipeff_1_w_lg_w_q_range931w932w & wire_y_pipeff_1_w_lg_w_q_range925w926w & wire_y_pipeff_1_w_lg_w_q_range919w920w & wire_y_pipeff_1_w_lg_w_q_range913w914w & wire_y_pipeff_1_w_lg_w_q_range907w908w & wire_y_pipeff_1_w_lg_w_q_range901w902w & wire_y_pipeff_1_w_lg_w_q_range895w896w & wire_y_pipeff_1_w_lg_w_q_range889w890w & wire_y_pipeff_1_w_lg_w_q_range883w884w & wire_y_pipeff_1_w_lg_w_q_range877w878w & wire_y_pipeff_1_w_lg_w_q_range871w872w);
	x_prenodetwo_3_w <= ( wire_y_pipeff_2_w_lg_w_q_range1697w1698w & wire_y_pipeff_2_w_lg_w_q_range1697w1698w & wire_y_pipeff_2_w_lg_w_q_range1697w1698w & wire_y_pipeff_2_w_lg_w_q_range1697w1698w & wire_y_pipeff_2_w_lg_w_q_range1697w1698w & wire_y_pipeff_2_w_lg_w_q_range1895w1896w & wire_y_pipeff_2_w_lg_w_q_range1889w1890w & wire_y_pipeff_2_w_lg_w_q_range1883w1884w & wire_y_pipeff_2_w_lg_w_q_range1877w1878w & wire_y_pipeff_2_w_lg_w_q_range1871w1872w & wire_y_pipeff_2_w_lg_w_q_range1865w1866w & wire_y_pipeff_2_w_lg_w_q_range1859w1860w & wire_y_pipeff_2_w_lg_w_q_range1853w1854w & wire_y_pipeff_2_w_lg_w_q_range1847w1848w & wire_y_pipeff_2_w_lg_w_q_range1841w1842w & wire_y_pipeff_2_w_lg_w_q_range1835w1836w & wire_y_pipeff_2_w_lg_w_q_range1829w1830w & wire_y_pipeff_2_w_lg_w_q_range1823w1824w & wire_y_pipeff_2_w_lg_w_q_range1817w1818w & wire_y_pipeff_2_w_lg_w_q_range1811w1812w & wire_y_pipeff_2_w_lg_w_q_range1805w1806w & wire_y_pipeff_2_w_lg_w_q_range1799w1800w & wire_y_pipeff_2_w_lg_w_q_range1793w1794w & wire_y_pipeff_2_w_lg_w_q_range1787w1788w & wire_y_pipeff_2_w_lg_w_q_range1781w1782w & wire_y_pipeff_2_w_lg_w_q_range1775w1776w & wire_y_pipeff_2_w_lg_w_q_range1769w1770w & wire_y_pipeff_2_w_lg_w_q_range1763w1764w & wire_y_pipeff_2_w_lg_w_q_range1757w1758w & wire_y_pipeff_2_w_lg_w_q_range1751w1752w & wire_y_pipeff_2_w_lg_w_q_range1745w1746w & wire_y_pipeff_2_w_lg_w_q_range1739w1740w & wire_y_pipeff_2_w_lg_w_q_range1733w1734w & wire_y_pipeff_2_w_lg_w_q_range1727w1728w);
	x_prenodetwo_4_w <= ( wire_y_pipeff_3_w_lg_w_q_range2544w2545w & wire_y_pipeff_3_w_lg_w_q_range2544w2545w & wire_y_pipeff_3_w_lg_w_q_range2544w2545w & wire_y_pipeff_3_w_lg_w_q_range2544w2545w & wire_y_pipeff_3_w_lg_w_q_range2544w2545w & wire_y_pipeff_3_w_lg_w_q_range2544w2545w & wire_y_pipeff_3_w_lg_w_q_range2740w2741w & wire_y_pipeff_3_w_lg_w_q_range2734w2735w & wire_y_pipeff_3_w_lg_w_q_range2728w2729w & wire_y_pipeff_3_w_lg_w_q_range2722w2723w & wire_y_pipeff_3_w_lg_w_q_range2716w2717w & wire_y_pipeff_3_w_lg_w_q_range2710w2711w & wire_y_pipeff_3_w_lg_w_q_range2704w2705w & wire_y_pipeff_3_w_lg_w_q_range2698w2699w & wire_y_pipeff_3_w_lg_w_q_range2692w2693w & wire_y_pipeff_3_w_lg_w_q_range2686w2687w & wire_y_pipeff_3_w_lg_w_q_range2680w2681w & wire_y_pipeff_3_w_lg_w_q_range2674w2675w & wire_y_pipeff_3_w_lg_w_q_range2668w2669w & wire_y_pipeff_3_w_lg_w_q_range2662w2663w & wire_y_pipeff_3_w_lg_w_q_range2656w2657w & wire_y_pipeff_3_w_lg_w_q_range2650w2651w & wire_y_pipeff_3_w_lg_w_q_range2644w2645w & wire_y_pipeff_3_w_lg_w_q_range2638w2639w & wire_y_pipeff_3_w_lg_w_q_range2632w2633w & wire_y_pipeff_3_w_lg_w_q_range2626w2627w & wire_y_pipeff_3_w_lg_w_q_range2620w2621w & wire_y_pipeff_3_w_lg_w_q_range2614w2615w & wire_y_pipeff_3_w_lg_w_q_range2608w2609w & wire_y_pipeff_3_w_lg_w_q_range2602w2603w & wire_y_pipeff_3_w_lg_w_q_range2596w2597w & wire_y_pipeff_3_w_lg_w_q_range2590w2591w & wire_y_pipeff_3_w_lg_w_q_range2584w2585w & wire_y_pipeff_3_w_lg_w_q_range2578w2579w);
	x_prenodetwo_5_w <= ( wire_y_pipeff_4_w_lg_w_q_range3386w3387w & wire_y_pipeff_4_w_lg_w_q_range3386w3387w & wire_y_pipeff_4_w_lg_w_q_range3386w3387w & wire_y_pipeff_4_w_lg_w_q_range3386w3387w & wire_y_pipeff_4_w_lg_w_q_range3386w3387w & wire_y_pipeff_4_w_lg_w_q_range3386w3387w & wire_y_pipeff_4_w_lg_w_q_range3386w3387w & wire_y_pipeff_4_w_lg_w_q_range3580w3581w & wire_y_pipeff_4_w_lg_w_q_range3574w3575w & wire_y_pipeff_4_w_lg_w_q_range3568w3569w & wire_y_pipeff_4_w_lg_w_q_range3562w3563w & wire_y_pipeff_4_w_lg_w_q_range3556w3557w & wire_y_pipeff_4_w_lg_w_q_range3550w3551w & wire_y_pipeff_4_w_lg_w_q_range3544w3545w & wire_y_pipeff_4_w_lg_w_q_range3538w3539w & wire_y_pipeff_4_w_lg_w_q_range3532w3533w & wire_y_pipeff_4_w_lg_w_q_range3526w3527w & wire_y_pipeff_4_w_lg_w_q_range3520w3521w & wire_y_pipeff_4_w_lg_w_q_range3514w3515w & wire_y_pipeff_4_w_lg_w_q_range3508w3509w & wire_y_pipeff_4_w_lg_w_q_range3502w3503w & wire_y_pipeff_4_w_lg_w_q_range3496w3497w & wire_y_pipeff_4_w_lg_w_q_range3490w3491w & wire_y_pipeff_4_w_lg_w_q_range3484w3485w & wire_y_pipeff_4_w_lg_w_q_range3478w3479w & wire_y_pipeff_4_w_lg_w_q_range3472w3473w & wire_y_pipeff_4_w_lg_w_q_range3466w3467w & wire_y_pipeff_4_w_lg_w_q_range3460w3461w & wire_y_pipeff_4_w_lg_w_q_range3454w3455w & wire_y_pipeff_4_w_lg_w_q_range3448w3449w & wire_y_pipeff_4_w_lg_w_q_range3442w3443w & wire_y_pipeff_4_w_lg_w_q_range3436w3437w & wire_y_pipeff_4_w_lg_w_q_range3430w3431w & wire_y_pipeff_4_w_lg_w_q_range3424w3425w);
	x_prenodetwo_6_w <= ( wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4223w4224w & wire_y_pipeff_5_w_lg_w_q_range4415w4416w & wire_y_pipeff_5_w_lg_w_q_range4409w4410w & wire_y_pipeff_5_w_lg_w_q_range4403w4404w & wire_y_pipeff_5_w_lg_w_q_range4397w4398w & wire_y_pipeff_5_w_lg_w_q_range4391w4392w & wire_y_pipeff_5_w_lg_w_q_range4385w4386w & wire_y_pipeff_5_w_lg_w_q_range4379w4380w & wire_y_pipeff_5_w_lg_w_q_range4373w4374w & wire_y_pipeff_5_w_lg_w_q_range4367w4368w & wire_y_pipeff_5_w_lg_w_q_range4361w4362w & wire_y_pipeff_5_w_lg_w_q_range4355w4356w & wire_y_pipeff_5_w_lg_w_q_range4349w4350w & wire_y_pipeff_5_w_lg_w_q_range4343w4344w & wire_y_pipeff_5_w_lg_w_q_range4337w4338w & wire_y_pipeff_5_w_lg_w_q_range4331w4332w & wire_y_pipeff_5_w_lg_w_q_range4325w4326w & wire_y_pipeff_5_w_lg_w_q_range4319w4320w & wire_y_pipeff_5_w_lg_w_q_range4313w4314w & wire_y_pipeff_5_w_lg_w_q_range4307w4308w & wire_y_pipeff_5_w_lg_w_q_range4301w4302w & wire_y_pipeff_5_w_lg_w_q_range4295w4296w & wire_y_pipeff_5_w_lg_w_q_range4289w4290w & wire_y_pipeff_5_w_lg_w_q_range4283w4284w & wire_y_pipeff_5_w_lg_w_q_range4277w4278w & wire_y_pipeff_5_w_lg_w_q_range4271w4272w & wire_y_pipeff_5_w_lg_w_q_range4265w4266w);
	x_prenodetwo_7_w <= ( wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5055w5056w & wire_y_pipeff_6_w_lg_w_q_range5245w5246w & wire_y_pipeff_6_w_lg_w_q_range5239w5240w & wire_y_pipeff_6_w_lg_w_q_range5233w5234w & wire_y_pipeff_6_w_lg_w_q_range5227w5228w & wire_y_pipeff_6_w_lg_w_q_range5221w5222w & wire_y_pipeff_6_w_lg_w_q_range5215w5216w & wire_y_pipeff_6_w_lg_w_q_range5209w5210w & wire_y_pipeff_6_w_lg_w_q_range5203w5204w & wire_y_pipeff_6_w_lg_w_q_range5197w5198w & wire_y_pipeff_6_w_lg_w_q_range5191w5192w & wire_y_pipeff_6_w_lg_w_q_range5185w5186w & wire_y_pipeff_6_w_lg_w_q_range5179w5180w & wire_y_pipeff_6_w_lg_w_q_range5173w5174w & wire_y_pipeff_6_w_lg_w_q_range5167w5168w & wire_y_pipeff_6_w_lg_w_q_range5161w5162w & wire_y_pipeff_6_w_lg_w_q_range5155w5156w & wire_y_pipeff_6_w_lg_w_q_range5149w5150w & wire_y_pipeff_6_w_lg_w_q_range5143w5144w & wire_y_pipeff_6_w_lg_w_q_range5137w5138w & wire_y_pipeff_6_w_lg_w_q_range5131w5132w & wire_y_pipeff_6_w_lg_w_q_range5125w5126w & wire_y_pipeff_6_w_lg_w_q_range5119w5120w & wire_y_pipeff_6_w_lg_w_q_range5113w5114w & wire_y_pipeff_6_w_lg_w_q_range5107w5108w & wire_y_pipeff_6_w_lg_w_q_range5101w5102w);
	x_prenodetwo_8_w <= ( wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range5882w5883w & wire_y_pipeff_7_w_lg_w_q_range6070w6071w & wire_y_pipeff_7_w_lg_w_q_range6064w6065w & wire_y_pipeff_7_w_lg_w_q_range6058w6059w & wire_y_pipeff_7_w_lg_w_q_range6052w6053w & wire_y_pipeff_7_w_lg_w_q_range6046w6047w & wire_y_pipeff_7_w_lg_w_q_range6040w6041w & wire_y_pipeff_7_w_lg_w_q_range6034w6035w & wire_y_pipeff_7_w_lg_w_q_range6028w6029w & wire_y_pipeff_7_w_lg_w_q_range6022w6023w & wire_y_pipeff_7_w_lg_w_q_range6016w6017w & wire_y_pipeff_7_w_lg_w_q_range6010w6011w & wire_y_pipeff_7_w_lg_w_q_range6004w6005w & wire_y_pipeff_7_w_lg_w_q_range5998w5999w & wire_y_pipeff_7_w_lg_w_q_range5992w5993w & wire_y_pipeff_7_w_lg_w_q_range5986w5987w & wire_y_pipeff_7_w_lg_w_q_range5980w5981w & wire_y_pipeff_7_w_lg_w_q_range5974w5975w & wire_y_pipeff_7_w_lg_w_q_range5968w5969w & wire_y_pipeff_7_w_lg_w_q_range5962w5963w & wire_y_pipeff_7_w_lg_w_q_range5956w5957w & wire_y_pipeff_7_w_lg_w_q_range5950w5951w & wire_y_pipeff_7_w_lg_w_q_range5944w5945w & wire_y_pipeff_7_w_lg_w_q_range5938w5939w & wire_y_pipeff_7_w_lg_w_q_range5932w5933w);
	x_prenodetwo_9_w <= ( wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6704w6705w & wire_y_pipeff_8_w_lg_w_q_range6890w6891w & wire_y_pipeff_8_w_lg_w_q_range6884w6885w & wire_y_pipeff_8_w_lg_w_q_range6878w6879w & wire_y_pipeff_8_w_lg_w_q_range6872w6873w & wire_y_pipeff_8_w_lg_w_q_range6866w6867w & wire_y_pipeff_8_w_lg_w_q_range6860w6861w & wire_y_pipeff_8_w_lg_w_q_range6854w6855w & wire_y_pipeff_8_w_lg_w_q_range6848w6849w & wire_y_pipeff_8_w_lg_w_q_range6842w6843w & wire_y_pipeff_8_w_lg_w_q_range6836w6837w & wire_y_pipeff_8_w_lg_w_q_range6830w6831w & wire_y_pipeff_8_w_lg_w_q_range6824w6825w & wire_y_pipeff_8_w_lg_w_q_range6818w6819w & wire_y_pipeff_8_w_lg_w_q_range6812w6813w & wire_y_pipeff_8_w_lg_w_q_range6806w6807w & wire_y_pipeff_8_w_lg_w_q_range6800w6801w & wire_y_pipeff_8_w_lg_w_q_range6794w6795w & wire_y_pipeff_8_w_lg_w_q_range6788w6789w & wire_y_pipeff_8_w_lg_w_q_range6782w6783w & wire_y_pipeff_8_w_lg_w_q_range6776w6777w & wire_y_pipeff_8_w_lg_w_q_range6770w6771w & wire_y_pipeff_8_w_lg_w_q_range6764w6765w & wire_y_pipeff_8_w_lg_w_q_range6758w6759w);
	x_start_node_w <= wire_cxs_value;
	x_subnode_10_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8052w8325w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8044w8317w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8036w8309w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8028w8301w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8020w8293w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8012w8285w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range8004w8277w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7996w8269w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7988w8261w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7980w8253w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7972w8245w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7964w8237w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7956w8229w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7948w8221w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7940w8213w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7932w8205w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7924w8197w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7916w8189w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7908w8181w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7900w8173w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7892w8165w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7884w8157w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7876w8149w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7868w8141w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7860w8133w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7852w8125w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7844w8117w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7836w8109w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7828w8101w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7820w8093w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7812w8085w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7804w8077w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7796w8069w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7786w8058w);
	x_subnode_11_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8859w9132w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8851w9124w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8843w9116w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8835w9108w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8827w9100w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8819w9092w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8811w9084w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8803w9076w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8795w9068w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8787w9060w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8779w9052w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8771w9044w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8763w9036w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8755w9028w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8747w9020w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8739w9012w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8731w9004w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8723w8996w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8715w8988w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8707w8980w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8699w8972w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8691w8964w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8683w8956w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8675w8948w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8667w8940w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8659w8932w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8651w8924w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8643w8916w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8635w8908w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8627w8900w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8619w8892w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8611w8884w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8603w8876w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8593w8865w);
	x_subnode_12_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9661w9934w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9653w9926w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9645w9918w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9637w9910w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9629w9902w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9621w9894w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9613w9886w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9605w9878w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9597w9870w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9589w9862w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9581w9854w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9573w9846w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9565w9838w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9557w9830w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9549w9822w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9541w9814w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9533w9806w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9525w9798w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9517w9790w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9509w9782w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9501w9774w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9493w9766w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9485w9758w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9477w9750w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9469w9742w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9461w9734w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9453w9726w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9445w9718w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9437w9710w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9429w9702w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9421w9694w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9413w9686w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9405w9678w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range9395w9667w);
	x_subnode_13_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10458w10731w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10450w10723w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10442w10715w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10434w10707w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10426w10699w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10418w10691w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10410w10683w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10402w10675w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10394w10667w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10386w10659w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10378w10651w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10370w10643w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10362w10635w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10354w10627w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10346w10619w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10338w10611w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10330w10603w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10322w10595w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10314w10587w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10306w10579w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10298w10571w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10290w10563w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10282w10555w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10274w10547w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10266w10539w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10258w10531w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10250w10523w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10242w10515w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10234w10507w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10226w10499w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10218w10491w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10210w10483w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10202w10475w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range10192w10464w
);
	x_subnode_2_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1416w1689w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1408w1681w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1400w1673w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1392w1665w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1384w1657w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1376w1649w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1368w1641w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1360w1633w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1352w1625w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1344w1617w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1336w1609w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1328w1601w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1320w1593w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1312w1585w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1304w1577w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1296w1569w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1288w1561w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1280w1553w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1272w1545w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1264w1537w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1256w1529w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1248w1521w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1240w1513w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1232w1505w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1224w1497w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1216w1489w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1208w1481w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1200w1473w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1192w1465w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1184w1457w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1176w1449w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1168w1441w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1160w1433w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1150w1422w);
	x_subnode_3_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2263w2536w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2255w2528w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2247w2520w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2239w2512w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2231w2504w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2223w2496w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2215w2488w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2207w2480w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2199w2472w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2191w2464w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2183w2456w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2175w2448w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2167w2440w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2159w2432w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2151w2424w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2143w2416w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2135w2408w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2127w2400w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2119w2392w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2111w2384w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2103w2376w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2095w2368w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2087w2360w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2079w2352w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2071w2344w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2063w2336w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2055w2328w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2047w2320w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2039w2312w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2031w2304w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2023w2296w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2015w2288w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2007w2280w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1997w2269w);
	x_subnode_4_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3105w3378w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3097w3370w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3089w3362w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3081w3354w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3073w3346w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3065w3338w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3057w3330w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3049w3322w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3041w3314w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3033w3306w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3025w3298w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3017w3290w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3009w3282w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range3001w3274w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2993w3266w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2985w3258w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2977w3250w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2969w3242w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2961w3234w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2953w3226w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2945w3218w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2937w3210w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2929w3202w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2921w3194w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2913w3186w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2905w3178w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2897w3170w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2889w3162w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2881w3154w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2873w3146w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2865w3138w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2857w3130w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2849w3122w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2839w3111w);
	x_subnode_5_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3942w4215w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3934w4207w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3926w4199w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3918w4191w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3910w4183w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3902w4175w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3894w4167w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3886w4159w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3878w4151w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3870w4143w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3862w4135w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3854w4127w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3846w4119w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3838w4111w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3830w4103w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3822w4095w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3814w4087w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3806w4079w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3798w4071w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3790w4063w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3782w4055w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3774w4047w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3766w4039w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3758w4031w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3750w4023w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3742w4015w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3734w4007w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3726w3999w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3718w3991w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3710w3983w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3702w3975w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3694w3967w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3686w3959w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3676w3948w);
	x_subnode_6_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4774w5047w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4766w5039w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4758w5031w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4750w5023w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4742w5015w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4734w5007w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4726w4999w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4718w4991w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4710w4983w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4702w4975w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4694w4967w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4686w4959w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4678w4951w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4670w4943w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4662w4935w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4654w4927w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4646w4919w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4638w4911w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4630w4903w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4622w4895w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4614w4887w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4606w4879w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4598w4871w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4590w4863w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4582w4855w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4574w4847w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4566w4839w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4558w4831w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4550w4823w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4542w4815w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4534w4807w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4526w4799w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4518w4791w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4508w4780w);
	x_subnode_7_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5601w5874w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5593w5866w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5585w5858w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5577w5850w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5569w5842w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5561w5834w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5553w5826w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5545w5818w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5537w5810w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5529w5802w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5521w5794w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5513w5786w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5505w5778w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5497w5770w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5489w5762w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5481w5754w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5473w5746w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5465w5738w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5457w5730w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5449w5722w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5441w5714w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5433w5706w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5425w5698w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5417w5690w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5409w5682w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5401w5674w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5393w5666w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5385w5658w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5377w5650w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5369w5642w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5361w5634w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5353w5626w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5345w5618w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5335w5607w);
	x_subnode_8_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6423w6696w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6415w6688w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6407w6680w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6399w6672w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6391w6664w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6383w6656w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6375w6648w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6367w6640w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6359w6632w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6351w6624w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6343w6616w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6335w6608w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6327w6600w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6319w6592w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6311w6584w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6303w6576w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6295w6568w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6287w6560w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6279w6552w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6271w6544w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6263w6536w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6255w6528w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6247w6520w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6239w6512w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6231w6504w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6223w6496w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6215w6488w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6207w6480w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6199w6472w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6191w6464w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6183w6456w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6175w6448w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6167w6440w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range6157w6429w);
	x_subnode_9_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7240w7513w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7232w7505w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7224w7497w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7216w7489w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7208w7481w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7200w7473w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7192w7465w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7184w7457w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7176w7449w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7168w7441w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7160w7433w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7152w7425w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7144w7417w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7136w7409w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7128w7401w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7120w7393w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7112w7385w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7104w7377w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7096w7369w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7088w7361w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7080w7353w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7072w7345w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7064w7337w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7056w7329w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7048w7321w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7040w7313w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7032w7305w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7024w7297w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7016w7289w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7008w7281w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range7000w7273w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6992w7265w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6984w7257w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6974w7246w);
	y_pipenode_10_w <= wire_y_pipenode_10_add_result;
	y_pipenode_11_w <= wire_y_pipenode_11_add_result;
	y_pipenode_12_w <= wire_y_pipenode_12_add_result;
	y_pipenode_13_w <= wire_y_pipenode_13_add_result;
	y_pipenode_2_w <= wire_y_pipenode_2_add_result;
	y_pipenode_3_w <= wire_y_pipenode_3_add_result;
	y_pipenode_4_w <= wire_y_pipenode_4_add_result;
	y_pipenode_5_w <= wire_y_pipenode_5_add_result;
	y_pipenode_6_w <= wire_y_pipenode_6_add_result;
	y_pipenode_7_w <= wire_y_pipenode_7_add_result;
	y_pipenode_8_w <= wire_y_pipenode_8_add_result;
	y_pipenode_9_w <= wire_y_pipenode_9_add_result;
	y_prenode_10_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7543w8054w8055w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7541w8046w8047w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7539w8038w8039w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7537w8030w8031w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7535w8022w8023w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7533w8014w8015w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7531w8006w8007w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7529w7998w7999w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7526w7990w7991w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7712w7982w7983w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7709w7974w7975w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7703w7966w7967w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7697w7958w7959w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7691w7950w7951w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7685w7942w7943w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7679w7934w7935w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7673w7926w7927w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7667w7918w7919w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7661w7910w7911w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7655w7902w7903w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7649w7894w7895w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7643w7886w7887w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7637w7878w7879w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7631w7870w7871w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7625w7862w7863w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7619w7854w7855w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7613w7846w7847w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7607w7838w7839w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7601w7830w7831w
 & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7595w7822w7823w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7589w7814w7815w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7583w7806w7807w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7577w7798w7799w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7572w7789w7790w);
	y_prenode_11_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8357w8861w8862w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8355w8853w8854w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8353w8845w8846w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8351w8837w8838w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8349w8829w8830w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8347w8821w8822w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8345w8813w8814w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8343w8805w8806w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8341w8797w8798w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8338w8789w8790w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8522w8781w8782w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8519w8773w8774w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8513w8765w8766w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8507w8757w8758w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8501w8749w8750w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8495w8741w8742w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8489w8733w8734w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8483w8725w8726w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8477w8717w8718w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8471w8709w8710w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8465w8701w8702w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8459w8693w8694w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8453w8685w8686w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8447w8677w8678w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8441w8669w8670w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8435w8661w8662w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8429w8653w8654w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8423w8645w8646w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8417w8637w8638w
 & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8411w8629w8630w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8405w8621w8622w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8399w8613w8614w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8393w8605w8606w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range8388w8596w8597w);
	y_prenode_12_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9166w9663w9664w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9164w9655w9656w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9162w9647w9648w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9160w9639w9640w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9158w9631w9632w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9156w9623w9624w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9154w9615w9616w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9152w9607w9608w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9150w9599w9600w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9148w9591w9592w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9145w9583w9584w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9327w9575w9576w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9324w9567w9568w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9318w9559w9560w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9312w9551w9552w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9306w9543w9544w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9300w9535w9536w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9294w9527w9528w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9288w9519w9520w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9282w9511w9512w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9276w9503w9504w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9270w9495w9496w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9264w9487w9488w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9258w9479w9480w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9252w9471w9472w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9246w9463w9464w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9240w9455w9456w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9234w9447w9448w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9228w9439w9440w
 & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9222w9431w9432w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9216w9423w9424w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9210w9415w9416w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9204w9407w9408w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range9199w9398w9399w);
	y_prenode_13_w <= ( wire_ccc_cordic_m_w10461w & wire_ccc_cordic_m_w10453w & wire_ccc_cordic_m_w10445w & wire_ccc_cordic_m_w10437w & wire_ccc_cordic_m_w10429w & wire_ccc_cordic_m_w10421w & wire_ccc_cordic_m_w10413w & wire_ccc_cordic_m_w10405w & wire_ccc_cordic_m_w10397w & wire_ccc_cordic_m_w10389w & wire_ccc_cordic_m_w10381w & wire_ccc_cordic_m_w10373w & wire_ccc_cordic_m_w10365w & wire_ccc_cordic_m_w10357w & wire_ccc_cordic_m_w10349w & wire_ccc_cordic_m_w10341w & wire_ccc_cordic_m_w10333w & wire_ccc_cordic_m_w10325w & wire_ccc_cordic_m_w10317w & wire_ccc_cordic_m_w10309w & wire_ccc_cordic_m_w10301w & wire_ccc_cordic_m_w10293w & wire_ccc_cordic_m_w10285w & wire_ccc_cordic_m_w10277w & wire_ccc_cordic_m_w10269w & wire_ccc_cordic_m_w10261w & wire_ccc_cordic_m_w10253w & wire_ccc_cordic_m_w10245w & wire_ccc_cordic_m_w10237w & wire_ccc_cordic_m_w10229w & wire_ccc_cordic_m_w10221w & wire_ccc_cordic_m_w10213w & wire_ccc_cordic_m_w10205w & wire_ccc_cordic_m_w10196w);
	y_prenode_2_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range850w1418w1419w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1052w1410w1411w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1049w1402w1403w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1043w1394w1395w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1037w1386w1387w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1031w1378w1379w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1025w1370w1371w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1019w1362w1363w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1013w1354w1355w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1007w1346w1347w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range1001w1338w1339w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range995w1330w1331w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range989w1322w1323w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range983w1314w1315w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range977w1306w1307w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range971w1298w1299w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range965w1290w1291w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range959w1282w1283w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range953w1274w1275w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range947w1266w1267w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range941w1258w1259w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range935w1250w1251w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range929w1242w1243w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range923w1234w1235w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range917w1226w1227w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range911w1218w1219w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range905w1210w1211w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range899w1202w1203w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range893w1194w1195w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range887w1186w1187w
 & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range881w1178w1179w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range875w1170w1171w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range869w1162w1163w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range864w1153w1154w);
	y_prenode_3_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1705w2265w2266w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1702w2257w2258w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1902w2249w2250w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1899w2241w2242w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1893w2233w2234w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1887w2225w2226w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1881w2217w2218w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1875w2209w2210w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1869w2201w2202w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1863w2193w2194w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1857w2185w2186w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1851w2177w2178w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1845w2169w2170w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1839w2161w2162w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1833w2153w2154w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1827w2145w2146w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1821w2137w2138w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1815w2129w2130w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1809w2121w2122w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1803w2113w2114w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1797w2105w2106w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1791w2097w2098w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1785w2089w2090w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1779w2081w2082w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1773w2073w2074w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1767w2065w2066w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1761w2057w2058w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1755w2049w2050w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1749w2041w2042w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1743w2033w2034w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1737w2025w2026w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1731w2017w2018w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1725w2009w2010w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1720w2000w2001w);
	y_prenode_4_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2554w3107w3108w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2552w3099w3100w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2549w3091w3092w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2747w3083w3084w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2744w3075w3076w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2738w3067w3068w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2732w3059w3060w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2726w3051w3052w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2720w3043w3044w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2714w3035w3036w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2708w3027w3028w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2702w3019w3020w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2696w3011w3012w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2690w3003w3004w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2684w2995w2996w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2678w2987w2988w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2672w2979w2980w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2666w2971w2972w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2660w2963w2964w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2654w2955w2956w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2648w2947w2948w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2642w2939w2940w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2636w2931w2932w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2630w2923w2924w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2624w2915w2916w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2618w2907w2908w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2612w2899w2900w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2606w2891w2892w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2600w2883w2884w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2594w2875w2876w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2588w2867w2868w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2582w2859w2860w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2576w2851w2852w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2571w2842w2843w);
	y_prenode_5_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3398w3944w3945w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3396w3936w3937w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3394w3928w3929w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3391w3920w3921w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3587w3912w3913w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3584w3904w3905w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3578w3896w3897w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3572w3888w3889w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3566w3880w3881w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3560w3872w3873w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3554w3864w3865w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3548w3856w3857w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3542w3848w3849w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3536w3840w3841w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3530w3832w3833w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3524w3824w3825w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3518w3816w3817w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3512w3808w3809w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3506w3800w3801w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3500w3792w3793w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3494w3784w3785w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3488w3776w3777w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3482w3768w3769w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3476w3760w3761w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3470w3752w3753w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3464w3744w3745w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3458w3736w3737w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3452w3728w3729w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3446w3720w3721w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3440w3712w3713w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3434w3704w3705w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3428w3696w3697w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3422w3688w3689w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3417w3679w3680w);
	y_prenode_6_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4237w4776w4777w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4235w4768w4769w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4233w4760w4761w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4231w4752w4753w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4228w4744w4745w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4422w4736w4737w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4419w4728w4729w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4413w4720w4721w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4407w4712w4713w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4401w4704w4705w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4395w4696w4697w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4389w4688w4689w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4383w4680w4681w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4377w4672w4673w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4371w4664w4665w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4365w4656w4657w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4359w4648w4649w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4353w4640w4641w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4347w4632w4633w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4341w4624w4625w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4335w4616w4617w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4329w4608w4609w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4323w4600w4601w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4317w4592w4593w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4311w4584w4585w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4305w4576w4577w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4299w4568w4569w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4293w4560w4561w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4287w4552w4553w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4281w4544w4545w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4275w4536w4537w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4269w4528w4529w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4263w4520w4521w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4258w4511w4512w);
	y_prenode_7_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5071w5603w5604w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5069w5595w5596w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5067w5587w5588w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5065w5579w5580w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5063w5571w5572w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5060w5563w5564w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5252w5555w5556w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5249w5547w5548w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5243w5539w5540w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5237w5531w5532w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5231w5523w5524w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5225w5515w5516w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5219w5507w5508w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5213w5499w5500w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5207w5491w5492w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5201w5483w5484w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5195w5475w5476w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5189w5467w5468w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5183w5459w5460w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5177w5451w5452w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5171w5443w5444w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5165w5435w5436w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5159w5427w5428w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5153w5419w5420w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5147w5411w5412w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5141w5403w5404w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5135w5395w5396w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5129w5387w5388w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5123w5379w5380w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5117w5371w5372w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5111w5363w5364w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5105w5355w5356w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5099w5347w5348w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range5094w5338w5339w);
	y_prenode_8_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5900w6425w6426w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5898w6417w6418w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5896w6409w6410w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5894w6401w6402w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5892w6393w6394w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5890w6385w6386w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5887w6377w6378w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6077w6369w6370w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6074w6361w6362w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6068w6353w6354w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6062w6345w6346w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6056w6337w6338w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6050w6329w6330w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6044w6321w6322w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6038w6313w6314w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6032w6305w6306w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6026w6297w6298w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6020w6289w6290w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6014w6281w6282w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6008w6273w6274w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range6002w6265w6266w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5996w6257w6258w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5990w6249w6250w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5984w6241w6242w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5978w6233w6234w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5972w6225w6226w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5966w6217w6218w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5960w6209w6210w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5954w6201w6202w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5948w6193w6194w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5942w6185w6186w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5936w6177w6178w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5930w6169w6170w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5925w6160w6161w);
	y_prenode_9_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6724w7242w7243w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6722w7234w7235w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6720w7226w7227w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6718w7218w7219w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6716w7210w7211w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6714w7202w7203w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6712w7194w7195w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6709w7186w7187w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6897w7178w7179w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6894w7170w7171w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6888w7162w7163w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6882w7154w7155w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6876w7146w7147w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6870w7138w7139w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6864w7130w7131w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6858w7122w7123w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6852w7114w7115w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6846w7106w7107w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6840w7098w7099w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6834w7090w7091w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6828w7082w7083w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6822w7074w7075w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6816w7066w7067w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6810w7058w7059w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6804w7050w7051w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6798w7042w7043w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6792w7034w7035w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6786w7026w7027w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6780w7018w7019w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6774w7010w7011w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6768w7002w7003w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6762w6994w6995w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6756w6986w6987w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6751w6977w6978w);
	y_prenodeone_10_w <= ( x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33 DOWNTO 9));
	y_prenodeone_11_w <= ( x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33 DOWNTO 10));
	y_prenodeone_12_w <= ( x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33 DOWNTO 11));
	y_prenodeone_13_w <= ( x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33 DOWNTO 12));
	y_prenodeone_2_w <= ( x_pipeff_1(33) & x_pipeff_1(33 DOWNTO 1));
	y_prenodeone_3_w <= ( x_pipeff_2(33) & x_pipeff_2(33) & x_pipeff_2(33 DOWNTO 2));
	y_prenodeone_4_w <= ( x_pipeff_3(33) & x_pipeff_3(33) & x_pipeff_3(33) & x_pipeff_3(33 DOWNTO 3));
	y_prenodeone_5_w <= ( x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33 DOWNTO 4));
	y_prenodeone_6_w <= ( x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33 DOWNTO 5));
	y_prenodeone_7_w <= ( x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33 DOWNTO 6));
	y_prenodeone_8_w <= ( x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33 DOWNTO 7));
	y_prenodeone_9_w <= ( x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33 DOWNTO 8));
	y_prenodetwo_10_w <= ( x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33) & x_pipeff_9(33 DOWNTO 11));
	y_prenodetwo_11_w <= ( x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33) & x_pipeff_10(33 DOWNTO 12));
	y_prenodetwo_12_w <= ( x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33) & x_pipeff_11(33 DOWNTO 13));
	y_prenodetwo_13_w <= ( x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33) & x_pipeff_12(33 DOWNTO 14));
	y_prenodetwo_2_w <= ( x_pipeff_1(33) & x_pipeff_1(33) & x_pipeff_1(33) & x_pipeff_1(33 DOWNTO 3));
	y_prenodetwo_3_w <= ( x_pipeff_2(33) & x_pipeff_2(33) & x_pipeff_2(33) & x_pipeff_2(33) & x_pipeff_2(33 DOWNTO 4));
	y_prenodetwo_4_w <= ( x_pipeff_3(33) & x_pipeff_3(33) & x_pipeff_3(33) & x_pipeff_3(33) & x_pipeff_3(33) & x_pipeff_3(33 DOWNTO 5));
	y_prenodetwo_5_w <= ( x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33) & x_pipeff_4(33 DOWNTO 6));
	y_prenodetwo_6_w <= ( x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33) & x_pipeff_5(33 DOWNTO 7));
	y_prenodetwo_7_w <= ( x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33) & x_pipeff_6(33 DOWNTO 8));
	y_prenodetwo_8_w <= ( x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33) & x_pipeff_7(33 DOWNTO 9));
	y_prenodetwo_9_w <= ( x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33) & x_pipeff_8(33 DOWNTO 10));
	y_subnode_10_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8056w8327w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8048w8319w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8040w8311w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8032w8303w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8024w8295w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8016w8287w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8008w8279w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range8000w8271w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7992w8263w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7984w8255w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7976w8247w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7968w8239w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7960w8231w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7952w8223w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7944w8215w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7936w8207w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7928w8199w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7920w8191w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7912w8183w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7904w8175w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7896w8167w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7888w8159w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7880w8151w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7872w8143w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7864w8135w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7856w8127w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7848w8119w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7840w8111w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7832w8103w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7824w8095w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7816w8087w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7808w8079w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7800w8071w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7791w8061w);
	y_subnode_11_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8863w9134w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8855w9126w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8847w9118w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8839w9110w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8831w9102w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8823w9094w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8815w9086w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8807w9078w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8799w9070w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8791w9062w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8783w9054w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8775w9046w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8767w9038w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8759w9030w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8751w9022w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8743w9014w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8735w9006w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8727w8998w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8719w8990w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8711w8982w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8703w8974w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8695w8966w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8687w8958w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8679w8950w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8671w8942w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8663w8934w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8655w8926w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8647w8918w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8639w8910w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8631w8902w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8623w8894w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8615w8886w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8607w8878w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8598w8868w);
	y_subnode_12_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9665w9936w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9657w9928w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9649w9920w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9641w9912w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9633w9904w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9625w9896w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9617w9888w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9609w9880w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9601w9872w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9593w9864w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9585w9856w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9577w9848w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9569w9840w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9561w9832w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9553w9824w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9545w9816w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9537w9808w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9529w9800w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9521w9792w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9513w9784w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9505w9776w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9497w9768w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9489w9760w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9481w9752w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9473w9744w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9465w9736w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9457w9728w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9449w9720w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9441w9712w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9433w9704w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9425w9696w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9417w9688w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9409w9680w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range9400w9670w);
	y_subnode_13_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10462w10733w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10454w10725w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10446w10717w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10438w10709w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10430w10701w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10422w10693w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10414w10685w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10406w10677w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10398w10669w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10390w10661w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10382w10653w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10374w10645w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10366w10637w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10358w10629w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10350w10621w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10342w10613w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10334w10605w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10326w10597w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10318w10589w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10310w10581w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10302w10573w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10294w10565w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10286w10557w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10278w10549w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10270w10541w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10262w10533w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10254w10525w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10246w10517w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10238w10509w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10230w10501w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10222w10493w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10214w10485w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10206w10477w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range10197w10467w
);
	y_subnode_1_w <= ( wire_x_pipeff_0_w_lg_w_q_range836w843w & wire_x_pipeff_0_w_lg_w_q_range831w841w & wire_x_pipeff_0_w_lg_w_lg_w_q_range826w838w839w & wire_x_pipeff_0_w_lg_w_lg_w_q_range821w833w834w & wire_x_pipeff_0_w_lg_w_lg_w_q_range816w828w829w & wire_x_pipeff_0_w_lg_w_lg_w_q_range811w823w824w & wire_x_pipeff_0_w_lg_w_lg_w_q_range806w818w819w & wire_x_pipeff_0_w_lg_w_lg_w_q_range801w813w814w & wire_x_pipeff_0_w_lg_w_lg_w_q_range796w808w809w & wire_x_pipeff_0_w_lg_w_lg_w_q_range791w803w804w & wire_x_pipeff_0_w_lg_w_lg_w_q_range786w798w799w & wire_x_pipeff_0_w_lg_w_lg_w_q_range781w793w794w & wire_x_pipeff_0_w_lg_w_lg_w_q_range776w788w789w & wire_x_pipeff_0_w_lg_w_lg_w_q_range771w783w784w & wire_x_pipeff_0_w_lg_w_lg_w_q_range766w778w779w & wire_x_pipeff_0_w_lg_w_lg_w_q_range761w773w774w & wire_x_pipeff_0_w_lg_w_lg_w_q_range756w768w769w & wire_x_pipeff_0_w_lg_w_lg_w_q_range751w763w764w & wire_x_pipeff_0_w_lg_w_lg_w_q_range746w758w759w & wire_x_pipeff_0_w_lg_w_lg_w_q_range741w753w754w & wire_x_pipeff_0_w_lg_w_lg_w_q_range736w748w749w & wire_x_pipeff_0_w_lg_w_lg_w_q_range731w743w744w & wire_x_pipeff_0_w_lg_w_lg_w_q_range726w738w739w & wire_x_pipeff_0_w_lg_w_lg_w_q_range721w733w734w & wire_x_pipeff_0_w_lg_w_lg_w_q_range716w728w729w & wire_x_pipeff_0_w_lg_w_lg_w_q_range711w723w724w & wire_x_pipeff_0_w_lg_w_lg_w_q_range706w718w719w & wire_x_pipeff_0_w_lg_w_lg_w_q_range701w713w714w & wire_x_pipeff_0_w_lg_w_lg_w_q_range696w708w709w & wire_x_pipeff_0_w_lg_w_lg_w_q_range691w703w704w & wire_x_pipeff_0_w_lg_w_lg_w_q_range685w698w699w & wire_x_pipeff_0_w_lg_w_lg_w_q_range677w693w694w & wire_x_pipeff_0_w_lg_w_lg_w_q_range687w688w689w & wire_x_pipeff_0_w_lg_w_lg_w_q_range680w681w682w);
	y_subnode_2_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1420w1691w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1412w1683w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1404w1675w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1396w1667w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1388w1659w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1380w1651w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1372w1643w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1364w1635w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1356w1627w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1348w1619w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1340w1611w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1332w1603w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1324w1595w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1316w1587w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1308w1579w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1300w1571w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1292w1563w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1284w1555w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1276w1547w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1268w1539w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1260w1531w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1252w1523w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1244w1515w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1236w1507w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1228w1499w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1220w1491w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1212w1483w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1204w1475w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1196w1467w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1188w1459w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1180w1451w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1172w1443w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1164w1435w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1155w1425w);
	y_subnode_3_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2267w2538w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2259w2530w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2251w2522w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2243w2514w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2235w2506w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2227w2498w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2219w2490w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2211w2482w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2203w2474w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2195w2466w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2187w2458w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2179w2450w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2171w2442w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2163w2434w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2155w2426w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2147w2418w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2139w2410w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2131w2402w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2123w2394w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2115w2386w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2107w2378w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2099w2370w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2091w2362w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2083w2354w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2075w2346w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2067w2338w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2059w2330w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2051w2322w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2043w2314w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2035w2306w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2027w2298w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2019w2290w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2011w2282w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2002w2272w);
	y_subnode_4_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3109w3380w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3101w3372w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3093w3364w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3085w3356w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3077w3348w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3069w3340w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3061w3332w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3053w3324w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3045w3316w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3037w3308w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3029w3300w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3021w3292w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3013w3284w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range3005w3276w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2997w3268w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2989w3260w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2981w3252w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2973w3244w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2965w3236w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2957w3228w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2949w3220w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2941w3212w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2933w3204w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2925w3196w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2917w3188w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2909w3180w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2901w3172w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2893w3164w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2885w3156w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2877w3148w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2869w3140w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2861w3132w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2853w3124w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2844w3114w);
	y_subnode_5_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3946w4217w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3938w4209w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3930w4201w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3922w4193w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3914w4185w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3906w4177w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3898w4169w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3890w4161w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3882w4153w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3874w4145w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3866w4137w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3858w4129w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3850w4121w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3842w4113w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3834w4105w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3826w4097w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3818w4089w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3810w4081w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3802w4073w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3794w4065w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3786w4057w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3778w4049w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3770w4041w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3762w4033w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3754w4025w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3746w4017w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3738w4009w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3730w4001w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3722w3993w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3714w3985w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3706w3977w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3698w3969w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3690w3961w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3681w3951w);
	y_subnode_6_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4778w5049w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4770w5041w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4762w5033w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4754w5025w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4746w5017w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4738w5009w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4730w5001w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4722w4993w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4714w4985w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4706w4977w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4698w4969w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4690w4961w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4682w4953w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4674w4945w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4666w4937w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4658w4929w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4650w4921w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4642w4913w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4634w4905w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4626w4897w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4618w4889w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4610w4881w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4602w4873w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4594w4865w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4586w4857w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4578w4849w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4570w4841w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4562w4833w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4554w4825w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4546w4817w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4538w4809w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4530w4801w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4522w4793w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4513w4783w);
	y_subnode_7_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5605w5876w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5597w5868w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5589w5860w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5581w5852w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5573w5844w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5565w5836w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5557w5828w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5549w5820w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5541w5812w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5533w5804w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5525w5796w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5517w5788w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5509w5780w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5501w5772w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5493w5764w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5485w5756w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5477w5748w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5469w5740w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5461w5732w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5453w5724w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5445w5716w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5437w5708w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5429w5700w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5421w5692w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5413w5684w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5405w5676w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5397w5668w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5389w5660w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5381w5652w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5373w5644w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5365w5636w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5357w5628w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5349w5620w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5340w5610w);
	y_subnode_8_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6427w6698w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6419w6690w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6411w6682w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6403w6674w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6395w6666w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6387w6658w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6379w6650w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6371w6642w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6363w6634w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6355w6626w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6347w6618w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6339w6610w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6331w6602w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6323w6594w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6315w6586w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6307w6578w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6299w6570w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6291w6562w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6283w6554w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6275w6546w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6267w6538w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6259w6530w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6251w6522w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6243w6514w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6235w6506w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6227w6498w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6219w6490w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6211w6482w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6203w6474w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6195w6466w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6187w6458w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6179w6450w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6171w6442w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range6162w6432w);
	y_subnode_9_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7244w7515w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7236w7507w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7228w7499w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7220w7491w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7212w7483w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7204w7475w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7196w7467w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7188w7459w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7180w7451w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7172w7443w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7164w7435w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7156w7427w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7148w7419w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7140w7411w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7132w7403w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7124w7395w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7116w7387w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7108w7379w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7100w7371w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7092w7363w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7084w7355w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7076w7347w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7068w7339w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7060w7331w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7052w7323w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7044w7315w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7036w7307w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7028w7299w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7020w7291w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7012w7283w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range7004w7275w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6996w7267w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6988w7259w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6979w7249w);
	z_pipenode_10_w <= wire_z_pipenode_10_add_result;
	z_pipenode_11_w <= wire_z_pipenode_11_add_result;
	z_pipenode_12_w <= wire_z_pipenode_12_add_result;
	z_pipenode_13_w <= wire_z_pipenode_13_add_result;
	z_pipenode_2_w <= wire_z_pipenode_2_add_result;
	z_pipenode_3_w <= wire_z_pipenode_3_add_result;
	z_pipenode_4_w <= wire_z_pipenode_4_add_result;
	z_pipenode_5_w <= wire_z_pipenode_5_add_result;
	z_pipenode_6_w <= wire_z_pipenode_6_add_result;
	z_pipenode_7_w <= wire_z_pipenode_7_add_result;
	z_pipenode_8_w <= wire_z_pipenode_8_add_result;
	z_pipenode_9_w <= wire_z_pipenode_9_add_result;
	z_subnode_10_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8329w8330w8331w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8321w8322w8323w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8313w8314w8315w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8305w8306w8307w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8297w8298w8299w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8289w8290w8291w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8281w8282w8283w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8273w8274w8275w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8265w8266w8267w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8257w8258w8259w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8249w8250w8251w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8241w8242w8243w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8233w8234w8235w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8225w8226w8227w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8217w8218w8219w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8209w8210w8211w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8201w8202w8203w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8193w8194w8195w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8185w8186w8187w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8177w8178w8179w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8169w8170w8171w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8161w8162w8163w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8153w8154w8155w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8145w8146w8147w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8137w8138w8139w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8129w8130w8131w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8121w8122w8123w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8113w8114w8115w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8105w8106w8107w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8097w8098w8099w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8089w8090w8091w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8081w8082w8083w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8073w8074w8075w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range8064w8065w8066w);
	z_subnode_11_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9136w9137w9138w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9128w9129w9130w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9120w9121w9122w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9112w9113w9114w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9104w9105w9106w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9096w9097w9098w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9088w9089w9090w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9080w9081w9082w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9072w9073w9074w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9064w9065w9066w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9056w9057w9058w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9048w9049w9050w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9040w9041w9042w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9032w9033w9034w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9024w9025w9026w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9016w9017w9018w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9008w9009w9010w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range9000w9001w9002w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8992w8993w8994w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8984w8985w8986w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8976w8977w8978w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8968w8969w8970w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8960w8961w8962w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8952w8953w8954w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8944w8945w8946w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8936w8937w8938w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8928w8929w8930w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8920w8921w8922w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8912w8913w8914w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8904w8905w8906w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8896w8897w8898w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8888w8889w8890w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8880w8881w8882w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8871w8872w8873w);
	z_subnode_12_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9938w9939w9940w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9930w9931w9932w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9922w9923w9924w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9914w9915w9916w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9906w9907w9908w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9898w9899w9900w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9890w9891w9892w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9882w9883w9884w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9874w9875w9876w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9866w9867w9868w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9858w9859w9860w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9850w9851w9852w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9842w9843w9844w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9834w9835w9836w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9826w9827w9828w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9818w9819w9820w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9810w9811w9812w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9802w9803w9804w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9794w9795w9796w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9786w9787w9788w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9778w9779w9780w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9770w9771w9772w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9762w9763w9764w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9754w9755w9756w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9746w9747w9748w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9738w9739w9740w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9730w9731w9732w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9722w9723w9724w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9714w9715w9716w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9706w9707w9708w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9698w9699w9700w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9690w9691w9692w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9682w9683w9684w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9673w9674w9675w);
	z_subnode_13_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10735w10736w10737w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10727w10728w10729w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10719w10720w10721w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10711w10712w10713w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10703w10704w10705w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10695w10696w10697w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10687w10688w10689w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10679w10680w10681w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10671w10672w10673w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10663w10664w10665w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10655w10656w10657w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10647w10648w10649w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10639w10640w10641w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10631w10632w10633w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10623w10624w10625w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10615w10616w10617w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10607w10608w10609w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10599w10600w10601w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10591w10592w10593w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10583w10584w10585w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10575w10576w10577w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10567w10568w10569w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10559w10560w10561w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10551w10552w10553w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10543w10544w10545w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10535w10536w10537w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10527w10528w10529w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10519w10520w10521w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10511w10512w10513w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10503w10504w10505w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10495w10496w10497w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10487w10488w10489w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10479w10480w10481w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range10470w10471w10472w);
	z_subnode_2_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1693w1694w1695w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1685w1686w1687w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1677w1678w1679w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1669w1670w1671w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1661w1662w1663w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1653w1654w1655w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1645w1646w1647w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1637w1638w1639w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1629w1630w1631w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1621w1622w1623w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1613w1614w1615w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1605w1606w1607w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1597w1598w1599w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1589w1590w1591w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1581w1582w1583w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1573w1574w1575w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1565w1566w1567w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1557w1558w1559w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1549w1550w1551w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1541w1542w1543w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1533w1534w1535w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1525w1526w1527w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1517w1518w1519w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1509w1510w1511w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1501w1502w1503w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1493w1494w1495w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1485w1486w1487w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1477w1478w1479w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1469w1470w1471w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1461w1462w1463w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1453w1454w1455w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1445w1446w1447w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1437w1438w1439w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1428w1429w1430w);
	z_subnode_3_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2540w2541w2542w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2532w2533w2534w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2524w2525w2526w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2516w2517w2518w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2508w2509w2510w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2500w2501w2502w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2492w2493w2494w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2484w2485w2486w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2476w2477w2478w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2468w2469w2470w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2460w2461w2462w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2452w2453w2454w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2444w2445w2446w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2436w2437w2438w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2428w2429w2430w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2420w2421w2422w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2412w2413w2414w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2404w2405w2406w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2396w2397w2398w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2388w2389w2390w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2380w2381w2382w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2372w2373w2374w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2364w2365w2366w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2356w2357w2358w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2348w2349w2350w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2340w2341w2342w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2332w2333w2334w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2324w2325w2326w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2316w2317w2318w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2308w2309w2310w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2300w2301w2302w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2292w2293w2294w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2284w2285w2286w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2275w2276w2277w);
	z_subnode_4_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3382w3383w3384w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3374w3375w3376w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3366w3367w3368w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3358w3359w3360w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3350w3351w3352w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3342w3343w3344w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3334w3335w3336w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3326w3327w3328w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3318w3319w3320w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3310w3311w3312w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3302w3303w3304w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3294w3295w3296w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3286w3287w3288w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3278w3279w3280w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3270w3271w3272w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3262w3263w3264w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3254w3255w3256w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3246w3247w3248w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3238w3239w3240w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3230w3231w3232w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3222w3223w3224w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3214w3215w3216w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3206w3207w3208w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3198w3199w3200w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3190w3191w3192w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3182w3183w3184w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3174w3175w3176w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3166w3167w3168w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3158w3159w3160w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3150w3151w3152w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3142w3143w3144w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3134w3135w3136w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3126w3127w3128w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3117w3118w3119w);
	z_subnode_5_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4219w4220w4221w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4211w4212w4213w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4203w4204w4205w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4195w4196w4197w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4187w4188w4189w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4179w4180w4181w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4171w4172w4173w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4163w4164w4165w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4155w4156w4157w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4147w4148w4149w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4139w4140w4141w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4131w4132w4133w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4123w4124w4125w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4115w4116w4117w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4107w4108w4109w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4099w4100w4101w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4091w4092w4093w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4083w4084w4085w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4075w4076w4077w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4067w4068w4069w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4059w4060w4061w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4051w4052w4053w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4043w4044w4045w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4035w4036w4037w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4027w4028w4029w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4019w4020w4021w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4011w4012w4013w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range4003w4004w4005w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3995w3996w3997w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3987w3988w3989w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3979w3980w3981w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3971w3972w3973w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3963w3964w3965w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3954w3955w3956w);
	z_subnode_6_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5051w5052w5053w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5043w5044w5045w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5035w5036w5037w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5027w5028w5029w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5019w5020w5021w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5011w5012w5013w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range5003w5004w5005w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4995w4996w4997w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4987w4988w4989w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4979w4980w4981w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4971w4972w4973w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4963w4964w4965w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4955w4956w4957w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4947w4948w4949w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4939w4940w4941w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4931w4932w4933w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4923w4924w4925w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4915w4916w4917w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4907w4908w4909w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4899w4900w4901w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4891w4892w4893w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4883w4884w4885w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4875w4876w4877w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4867w4868w4869w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4859w4860w4861w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4851w4852w4853w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4843w4844w4845w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4835w4836w4837w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4827w4828w4829w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4819w4820w4821w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4811w4812w4813w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4803w4804w4805w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4795w4796w4797w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4786w4787w4788w);
	z_subnode_7_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5878w5879w5880w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5870w5871w5872w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5862w5863w5864w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5854w5855w5856w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5846w5847w5848w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5838w5839w5840w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5830w5831w5832w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5822w5823w5824w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5814w5815w5816w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5806w5807w5808w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5798w5799w5800w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5790w5791w5792w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5782w5783w5784w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5774w5775w5776w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5766w5767w5768w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5758w5759w5760w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5750w5751w5752w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5742w5743w5744w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5734w5735w5736w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5726w5727w5728w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5718w5719w5720w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5710w5711w5712w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5702w5703w5704w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5694w5695w5696w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5686w5687w5688w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5678w5679w5680w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5670w5671w5672w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5662w5663w5664w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5654w5655w5656w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5646w5647w5648w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5638w5639w5640w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5630w5631w5632w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5622w5623w5624w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5613w5614w5615w);
	z_subnode_8_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6700w6701w6702w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6692w6693w6694w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6684w6685w6686w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6676w6677w6678w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6668w6669w6670w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6660w6661w6662w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6652w6653w6654w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6644w6645w6646w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6636w6637w6638w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6628w6629w6630w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6620w6621w6622w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6612w6613w6614w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6604w6605w6606w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6596w6597w6598w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6588w6589w6590w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6580w6581w6582w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6572w6573w6574w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6564w6565w6566w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6556w6557w6558w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6548w6549w6550w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6540w6541w6542w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6532w6533w6534w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6524w6525w6526w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6516w6517w6518w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6508w6509w6510w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6500w6501w6502w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6492w6493w6494w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6484w6485w6486w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6476w6477w6478w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6468w6469w6470w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6460w6461w6462w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6452w6453w6454w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6444w6445w6446w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6435w6436w6437w);
	z_subnode_9_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7517w7518w7519w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7509w7510w7511w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7501w7502w7503w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7493w7494w7495w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7485w7486w7487w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7477w7478w7479w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7469w7470w7471w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7461w7462w7463w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7453w7454w7455w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7445w7446w7447w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7437w7438w7439w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7429w7430w7431w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7421w7422w7423w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7413w7414w7415w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7405w7406w7407w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7397w7398w7399w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7389w7390w7391w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7381w7382w7383w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7373w7374w7375w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7365w7366w7367w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7357w7358w7359w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7349w7350w7351w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7341w7342w7343w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7333w7334w7335w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7325w7326w7327w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7317w7318w7319w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7309w7310w7311w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7301w7302w7303w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7293w7294w7295w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7285w7286w7287w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7277w7278w7279w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7269w7270w7271w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7261w7262w7263w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range7252w7253w7254w);
	wire_ccc_cordic_m_w_atannode_10_w_range8871w(0) <= atannode_10_w(0);
	wire_ccc_cordic_m_w_atannode_10_w_range8952w(0) <= atannode_10_w(10);
	wire_ccc_cordic_m_w_atannode_10_w_range8960w(0) <= atannode_10_w(11);
	wire_ccc_cordic_m_w_atannode_10_w_range8968w(0) <= atannode_10_w(12);
	wire_ccc_cordic_m_w_atannode_10_w_range8976w(0) <= atannode_10_w(13);
	wire_ccc_cordic_m_w_atannode_10_w_range8984w(0) <= atannode_10_w(14);
	wire_ccc_cordic_m_w_atannode_10_w_range8992w(0) <= atannode_10_w(15);
	wire_ccc_cordic_m_w_atannode_10_w_range9000w(0) <= atannode_10_w(16);
	wire_ccc_cordic_m_w_atannode_10_w_range9008w(0) <= atannode_10_w(17);
	wire_ccc_cordic_m_w_atannode_10_w_range9016w(0) <= atannode_10_w(18);
	wire_ccc_cordic_m_w_atannode_10_w_range9024w(0) <= atannode_10_w(19);
	wire_ccc_cordic_m_w_atannode_10_w_range8880w(0) <= atannode_10_w(1);
	wire_ccc_cordic_m_w_atannode_10_w_range9032w(0) <= atannode_10_w(20);
	wire_ccc_cordic_m_w_atannode_10_w_range9040w(0) <= atannode_10_w(21);
	wire_ccc_cordic_m_w_atannode_10_w_range9048w(0) <= atannode_10_w(22);
	wire_ccc_cordic_m_w_atannode_10_w_range9056w(0) <= atannode_10_w(23);
	wire_ccc_cordic_m_w_atannode_10_w_range9064w(0) <= atannode_10_w(24);
	wire_ccc_cordic_m_w_atannode_10_w_range9072w(0) <= atannode_10_w(25);
	wire_ccc_cordic_m_w_atannode_10_w_range9080w(0) <= atannode_10_w(26);
	wire_ccc_cordic_m_w_atannode_10_w_range9088w(0) <= atannode_10_w(27);
	wire_ccc_cordic_m_w_atannode_10_w_range9096w(0) <= atannode_10_w(28);
	wire_ccc_cordic_m_w_atannode_10_w_range9104w(0) <= atannode_10_w(29);
	wire_ccc_cordic_m_w_atannode_10_w_range8888w(0) <= atannode_10_w(2);
	wire_ccc_cordic_m_w_atannode_10_w_range9112w(0) <= atannode_10_w(30);
	wire_ccc_cordic_m_w_atannode_10_w_range9120w(0) <= atannode_10_w(31);
	wire_ccc_cordic_m_w_atannode_10_w_range9128w(0) <= atannode_10_w(32);
	wire_ccc_cordic_m_w_atannode_10_w_range9136w(0) <= atannode_10_w(33);
	wire_ccc_cordic_m_w_atannode_10_w_range8896w(0) <= atannode_10_w(3);
	wire_ccc_cordic_m_w_atannode_10_w_range8904w(0) <= atannode_10_w(4);
	wire_ccc_cordic_m_w_atannode_10_w_range8912w(0) <= atannode_10_w(5);
	wire_ccc_cordic_m_w_atannode_10_w_range8920w(0) <= atannode_10_w(6);
	wire_ccc_cordic_m_w_atannode_10_w_range8928w(0) <= atannode_10_w(7);
	wire_ccc_cordic_m_w_atannode_10_w_range8936w(0) <= atannode_10_w(8);
	wire_ccc_cordic_m_w_atannode_10_w_range8944w(0) <= atannode_10_w(9);
	wire_ccc_cordic_m_w_atannode_11_w_range9673w(0) <= atannode_11_w(0);
	wire_ccc_cordic_m_w_atannode_11_w_range9754w(0) <= atannode_11_w(10);
	wire_ccc_cordic_m_w_atannode_11_w_range9762w(0) <= atannode_11_w(11);
	wire_ccc_cordic_m_w_atannode_11_w_range9770w(0) <= atannode_11_w(12);
	wire_ccc_cordic_m_w_atannode_11_w_range9778w(0) <= atannode_11_w(13);
	wire_ccc_cordic_m_w_atannode_11_w_range9786w(0) <= atannode_11_w(14);
	wire_ccc_cordic_m_w_atannode_11_w_range9794w(0) <= atannode_11_w(15);
	wire_ccc_cordic_m_w_atannode_11_w_range9802w(0) <= atannode_11_w(16);
	wire_ccc_cordic_m_w_atannode_11_w_range9810w(0) <= atannode_11_w(17);
	wire_ccc_cordic_m_w_atannode_11_w_range9818w(0) <= atannode_11_w(18);
	wire_ccc_cordic_m_w_atannode_11_w_range9826w(0) <= atannode_11_w(19);
	wire_ccc_cordic_m_w_atannode_11_w_range9682w(0) <= atannode_11_w(1);
	wire_ccc_cordic_m_w_atannode_11_w_range9834w(0) <= atannode_11_w(20);
	wire_ccc_cordic_m_w_atannode_11_w_range9842w(0) <= atannode_11_w(21);
	wire_ccc_cordic_m_w_atannode_11_w_range9850w(0) <= atannode_11_w(22);
	wire_ccc_cordic_m_w_atannode_11_w_range9858w(0) <= atannode_11_w(23);
	wire_ccc_cordic_m_w_atannode_11_w_range9866w(0) <= atannode_11_w(24);
	wire_ccc_cordic_m_w_atannode_11_w_range9874w(0) <= atannode_11_w(25);
	wire_ccc_cordic_m_w_atannode_11_w_range9882w(0) <= atannode_11_w(26);
	wire_ccc_cordic_m_w_atannode_11_w_range9890w(0) <= atannode_11_w(27);
	wire_ccc_cordic_m_w_atannode_11_w_range9898w(0) <= atannode_11_w(28);
	wire_ccc_cordic_m_w_atannode_11_w_range9906w(0) <= atannode_11_w(29);
	wire_ccc_cordic_m_w_atannode_11_w_range9690w(0) <= atannode_11_w(2);
	wire_ccc_cordic_m_w_atannode_11_w_range9914w(0) <= atannode_11_w(30);
	wire_ccc_cordic_m_w_atannode_11_w_range9922w(0) <= atannode_11_w(31);
	wire_ccc_cordic_m_w_atannode_11_w_range9930w(0) <= atannode_11_w(32);
	wire_ccc_cordic_m_w_atannode_11_w_range9938w(0) <= atannode_11_w(33);
	wire_ccc_cordic_m_w_atannode_11_w_range9698w(0) <= atannode_11_w(3);
	wire_ccc_cordic_m_w_atannode_11_w_range9706w(0) <= atannode_11_w(4);
	wire_ccc_cordic_m_w_atannode_11_w_range9714w(0) <= atannode_11_w(5);
	wire_ccc_cordic_m_w_atannode_11_w_range9722w(0) <= atannode_11_w(6);
	wire_ccc_cordic_m_w_atannode_11_w_range9730w(0) <= atannode_11_w(7);
	wire_ccc_cordic_m_w_atannode_11_w_range9738w(0) <= atannode_11_w(8);
	wire_ccc_cordic_m_w_atannode_11_w_range9746w(0) <= atannode_11_w(9);
	wire_ccc_cordic_m_w_atannode_12_w_range10470w(0) <= atannode_12_w(0);
	wire_ccc_cordic_m_w_atannode_12_w_range10551w(0) <= atannode_12_w(10);
	wire_ccc_cordic_m_w_atannode_12_w_range10559w(0) <= atannode_12_w(11);
	wire_ccc_cordic_m_w_atannode_12_w_range10567w(0) <= atannode_12_w(12);
	wire_ccc_cordic_m_w_atannode_12_w_range10575w(0) <= atannode_12_w(13);
	wire_ccc_cordic_m_w_atannode_12_w_range10583w(0) <= atannode_12_w(14);
	wire_ccc_cordic_m_w_atannode_12_w_range10591w(0) <= atannode_12_w(15);
	wire_ccc_cordic_m_w_atannode_12_w_range10599w(0) <= atannode_12_w(16);
	wire_ccc_cordic_m_w_atannode_12_w_range10607w(0) <= atannode_12_w(17);
	wire_ccc_cordic_m_w_atannode_12_w_range10615w(0) <= atannode_12_w(18);
	wire_ccc_cordic_m_w_atannode_12_w_range10623w(0) <= atannode_12_w(19);
	wire_ccc_cordic_m_w_atannode_12_w_range10479w(0) <= atannode_12_w(1);
	wire_ccc_cordic_m_w_atannode_12_w_range10631w(0) <= atannode_12_w(20);
	wire_ccc_cordic_m_w_atannode_12_w_range10639w(0) <= atannode_12_w(21);
	wire_ccc_cordic_m_w_atannode_12_w_range10647w(0) <= atannode_12_w(22);
	wire_ccc_cordic_m_w_atannode_12_w_range10655w(0) <= atannode_12_w(23);
	wire_ccc_cordic_m_w_atannode_12_w_range10663w(0) <= atannode_12_w(24);
	wire_ccc_cordic_m_w_atannode_12_w_range10671w(0) <= atannode_12_w(25);
	wire_ccc_cordic_m_w_atannode_12_w_range10679w(0) <= atannode_12_w(26);
	wire_ccc_cordic_m_w_atannode_12_w_range10687w(0) <= atannode_12_w(27);
	wire_ccc_cordic_m_w_atannode_12_w_range10695w(0) <= atannode_12_w(28);
	wire_ccc_cordic_m_w_atannode_12_w_range10703w(0) <= atannode_12_w(29);
	wire_ccc_cordic_m_w_atannode_12_w_range10487w(0) <= atannode_12_w(2);
	wire_ccc_cordic_m_w_atannode_12_w_range10711w(0) <= atannode_12_w(30);
	wire_ccc_cordic_m_w_atannode_12_w_range10719w(0) <= atannode_12_w(31);
	wire_ccc_cordic_m_w_atannode_12_w_range10727w(0) <= atannode_12_w(32);
	wire_ccc_cordic_m_w_atannode_12_w_range10735w(0) <= atannode_12_w(33);
	wire_ccc_cordic_m_w_atannode_12_w_range10495w(0) <= atannode_12_w(3);
	wire_ccc_cordic_m_w_atannode_12_w_range10503w(0) <= atannode_12_w(4);
	wire_ccc_cordic_m_w_atannode_12_w_range10511w(0) <= atannode_12_w(5);
	wire_ccc_cordic_m_w_atannode_12_w_range10519w(0) <= atannode_12_w(6);
	wire_ccc_cordic_m_w_atannode_12_w_range10527w(0) <= atannode_12_w(7);
	wire_ccc_cordic_m_w_atannode_12_w_range10535w(0) <= atannode_12_w(8);
	wire_ccc_cordic_m_w_atannode_12_w_range10543w(0) <= atannode_12_w(9);
	wire_ccc_cordic_m_w_atannode_1_w_range1428w(0) <= atannode_1_w(0);
	wire_ccc_cordic_m_w_atannode_1_w_range1509w(0) <= atannode_1_w(10);
	wire_ccc_cordic_m_w_atannode_1_w_range1517w(0) <= atannode_1_w(11);
	wire_ccc_cordic_m_w_atannode_1_w_range1525w(0) <= atannode_1_w(12);
	wire_ccc_cordic_m_w_atannode_1_w_range1533w(0) <= atannode_1_w(13);
	wire_ccc_cordic_m_w_atannode_1_w_range1541w(0) <= atannode_1_w(14);
	wire_ccc_cordic_m_w_atannode_1_w_range1549w(0) <= atannode_1_w(15);
	wire_ccc_cordic_m_w_atannode_1_w_range1557w(0) <= atannode_1_w(16);
	wire_ccc_cordic_m_w_atannode_1_w_range1565w(0) <= atannode_1_w(17);
	wire_ccc_cordic_m_w_atannode_1_w_range1573w(0) <= atannode_1_w(18);
	wire_ccc_cordic_m_w_atannode_1_w_range1581w(0) <= atannode_1_w(19);
	wire_ccc_cordic_m_w_atannode_1_w_range1437w(0) <= atannode_1_w(1);
	wire_ccc_cordic_m_w_atannode_1_w_range1589w(0) <= atannode_1_w(20);
	wire_ccc_cordic_m_w_atannode_1_w_range1597w(0) <= atannode_1_w(21);
	wire_ccc_cordic_m_w_atannode_1_w_range1605w(0) <= atannode_1_w(22);
	wire_ccc_cordic_m_w_atannode_1_w_range1613w(0) <= atannode_1_w(23);
	wire_ccc_cordic_m_w_atannode_1_w_range1621w(0) <= atannode_1_w(24);
	wire_ccc_cordic_m_w_atannode_1_w_range1629w(0) <= atannode_1_w(25);
	wire_ccc_cordic_m_w_atannode_1_w_range1637w(0) <= atannode_1_w(26);
	wire_ccc_cordic_m_w_atannode_1_w_range1645w(0) <= atannode_1_w(27);
	wire_ccc_cordic_m_w_atannode_1_w_range1653w(0) <= atannode_1_w(28);
	wire_ccc_cordic_m_w_atannode_1_w_range1661w(0) <= atannode_1_w(29);
	wire_ccc_cordic_m_w_atannode_1_w_range1445w(0) <= atannode_1_w(2);
	wire_ccc_cordic_m_w_atannode_1_w_range1669w(0) <= atannode_1_w(30);
	wire_ccc_cordic_m_w_atannode_1_w_range1677w(0) <= atannode_1_w(31);
	wire_ccc_cordic_m_w_atannode_1_w_range1685w(0) <= atannode_1_w(32);
	wire_ccc_cordic_m_w_atannode_1_w_range1693w(0) <= atannode_1_w(33);
	wire_ccc_cordic_m_w_atannode_1_w_range1453w(0) <= atannode_1_w(3);
	wire_ccc_cordic_m_w_atannode_1_w_range1461w(0) <= atannode_1_w(4);
	wire_ccc_cordic_m_w_atannode_1_w_range1469w(0) <= atannode_1_w(5);
	wire_ccc_cordic_m_w_atannode_1_w_range1477w(0) <= atannode_1_w(6);
	wire_ccc_cordic_m_w_atannode_1_w_range1485w(0) <= atannode_1_w(7);
	wire_ccc_cordic_m_w_atannode_1_w_range1493w(0) <= atannode_1_w(8);
	wire_ccc_cordic_m_w_atannode_1_w_range1501w(0) <= atannode_1_w(9);
	wire_ccc_cordic_m_w_atannode_2_w_range2275w(0) <= atannode_2_w(0);
	wire_ccc_cordic_m_w_atannode_2_w_range2356w(0) <= atannode_2_w(10);
	wire_ccc_cordic_m_w_atannode_2_w_range2364w(0) <= atannode_2_w(11);
	wire_ccc_cordic_m_w_atannode_2_w_range2372w(0) <= atannode_2_w(12);
	wire_ccc_cordic_m_w_atannode_2_w_range2380w(0) <= atannode_2_w(13);
	wire_ccc_cordic_m_w_atannode_2_w_range2388w(0) <= atannode_2_w(14);
	wire_ccc_cordic_m_w_atannode_2_w_range2396w(0) <= atannode_2_w(15);
	wire_ccc_cordic_m_w_atannode_2_w_range2404w(0) <= atannode_2_w(16);
	wire_ccc_cordic_m_w_atannode_2_w_range2412w(0) <= atannode_2_w(17);
	wire_ccc_cordic_m_w_atannode_2_w_range2420w(0) <= atannode_2_w(18);
	wire_ccc_cordic_m_w_atannode_2_w_range2428w(0) <= atannode_2_w(19);
	wire_ccc_cordic_m_w_atannode_2_w_range2284w(0) <= atannode_2_w(1);
	wire_ccc_cordic_m_w_atannode_2_w_range2436w(0) <= atannode_2_w(20);
	wire_ccc_cordic_m_w_atannode_2_w_range2444w(0) <= atannode_2_w(21);
	wire_ccc_cordic_m_w_atannode_2_w_range2452w(0) <= atannode_2_w(22);
	wire_ccc_cordic_m_w_atannode_2_w_range2460w(0) <= atannode_2_w(23);
	wire_ccc_cordic_m_w_atannode_2_w_range2468w(0) <= atannode_2_w(24);
	wire_ccc_cordic_m_w_atannode_2_w_range2476w(0) <= atannode_2_w(25);
	wire_ccc_cordic_m_w_atannode_2_w_range2484w(0) <= atannode_2_w(26);
	wire_ccc_cordic_m_w_atannode_2_w_range2492w(0) <= atannode_2_w(27);
	wire_ccc_cordic_m_w_atannode_2_w_range2500w(0) <= atannode_2_w(28);
	wire_ccc_cordic_m_w_atannode_2_w_range2508w(0) <= atannode_2_w(29);
	wire_ccc_cordic_m_w_atannode_2_w_range2292w(0) <= atannode_2_w(2);
	wire_ccc_cordic_m_w_atannode_2_w_range2516w(0) <= atannode_2_w(30);
	wire_ccc_cordic_m_w_atannode_2_w_range2524w(0) <= atannode_2_w(31);
	wire_ccc_cordic_m_w_atannode_2_w_range2532w(0) <= atannode_2_w(32);
	wire_ccc_cordic_m_w_atannode_2_w_range2540w(0) <= atannode_2_w(33);
	wire_ccc_cordic_m_w_atannode_2_w_range2300w(0) <= atannode_2_w(3);
	wire_ccc_cordic_m_w_atannode_2_w_range2308w(0) <= atannode_2_w(4);
	wire_ccc_cordic_m_w_atannode_2_w_range2316w(0) <= atannode_2_w(5);
	wire_ccc_cordic_m_w_atannode_2_w_range2324w(0) <= atannode_2_w(6);
	wire_ccc_cordic_m_w_atannode_2_w_range2332w(0) <= atannode_2_w(7);
	wire_ccc_cordic_m_w_atannode_2_w_range2340w(0) <= atannode_2_w(8);
	wire_ccc_cordic_m_w_atannode_2_w_range2348w(0) <= atannode_2_w(9);
	wire_ccc_cordic_m_w_atannode_3_w_range3117w(0) <= atannode_3_w(0);
	wire_ccc_cordic_m_w_atannode_3_w_range3198w(0) <= atannode_3_w(10);
	wire_ccc_cordic_m_w_atannode_3_w_range3206w(0) <= atannode_3_w(11);
	wire_ccc_cordic_m_w_atannode_3_w_range3214w(0) <= atannode_3_w(12);
	wire_ccc_cordic_m_w_atannode_3_w_range3222w(0) <= atannode_3_w(13);
	wire_ccc_cordic_m_w_atannode_3_w_range3230w(0) <= atannode_3_w(14);
	wire_ccc_cordic_m_w_atannode_3_w_range3238w(0) <= atannode_3_w(15);
	wire_ccc_cordic_m_w_atannode_3_w_range3246w(0) <= atannode_3_w(16);
	wire_ccc_cordic_m_w_atannode_3_w_range3254w(0) <= atannode_3_w(17);
	wire_ccc_cordic_m_w_atannode_3_w_range3262w(0) <= atannode_3_w(18);
	wire_ccc_cordic_m_w_atannode_3_w_range3270w(0) <= atannode_3_w(19);
	wire_ccc_cordic_m_w_atannode_3_w_range3126w(0) <= atannode_3_w(1);
	wire_ccc_cordic_m_w_atannode_3_w_range3278w(0) <= atannode_3_w(20);
	wire_ccc_cordic_m_w_atannode_3_w_range3286w(0) <= atannode_3_w(21);
	wire_ccc_cordic_m_w_atannode_3_w_range3294w(0) <= atannode_3_w(22);
	wire_ccc_cordic_m_w_atannode_3_w_range3302w(0) <= atannode_3_w(23);
	wire_ccc_cordic_m_w_atannode_3_w_range3310w(0) <= atannode_3_w(24);
	wire_ccc_cordic_m_w_atannode_3_w_range3318w(0) <= atannode_3_w(25);
	wire_ccc_cordic_m_w_atannode_3_w_range3326w(0) <= atannode_3_w(26);
	wire_ccc_cordic_m_w_atannode_3_w_range3334w(0) <= atannode_3_w(27);
	wire_ccc_cordic_m_w_atannode_3_w_range3342w(0) <= atannode_3_w(28);
	wire_ccc_cordic_m_w_atannode_3_w_range3350w(0) <= atannode_3_w(29);
	wire_ccc_cordic_m_w_atannode_3_w_range3134w(0) <= atannode_3_w(2);
	wire_ccc_cordic_m_w_atannode_3_w_range3358w(0) <= atannode_3_w(30);
	wire_ccc_cordic_m_w_atannode_3_w_range3366w(0) <= atannode_3_w(31);
	wire_ccc_cordic_m_w_atannode_3_w_range3374w(0) <= atannode_3_w(32);
	wire_ccc_cordic_m_w_atannode_3_w_range3382w(0) <= atannode_3_w(33);
	wire_ccc_cordic_m_w_atannode_3_w_range3142w(0) <= atannode_3_w(3);
	wire_ccc_cordic_m_w_atannode_3_w_range3150w(0) <= atannode_3_w(4);
	wire_ccc_cordic_m_w_atannode_3_w_range3158w(0) <= atannode_3_w(5);
	wire_ccc_cordic_m_w_atannode_3_w_range3166w(0) <= atannode_3_w(6);
	wire_ccc_cordic_m_w_atannode_3_w_range3174w(0) <= atannode_3_w(7);
	wire_ccc_cordic_m_w_atannode_3_w_range3182w(0) <= atannode_3_w(8);
	wire_ccc_cordic_m_w_atannode_3_w_range3190w(0) <= atannode_3_w(9);
	wire_ccc_cordic_m_w_atannode_4_w_range3954w(0) <= atannode_4_w(0);
	wire_ccc_cordic_m_w_atannode_4_w_range4035w(0) <= atannode_4_w(10);
	wire_ccc_cordic_m_w_atannode_4_w_range4043w(0) <= atannode_4_w(11);
	wire_ccc_cordic_m_w_atannode_4_w_range4051w(0) <= atannode_4_w(12);
	wire_ccc_cordic_m_w_atannode_4_w_range4059w(0) <= atannode_4_w(13);
	wire_ccc_cordic_m_w_atannode_4_w_range4067w(0) <= atannode_4_w(14);
	wire_ccc_cordic_m_w_atannode_4_w_range4075w(0) <= atannode_4_w(15);
	wire_ccc_cordic_m_w_atannode_4_w_range4083w(0) <= atannode_4_w(16);
	wire_ccc_cordic_m_w_atannode_4_w_range4091w(0) <= atannode_4_w(17);
	wire_ccc_cordic_m_w_atannode_4_w_range4099w(0) <= atannode_4_w(18);
	wire_ccc_cordic_m_w_atannode_4_w_range4107w(0) <= atannode_4_w(19);
	wire_ccc_cordic_m_w_atannode_4_w_range3963w(0) <= atannode_4_w(1);
	wire_ccc_cordic_m_w_atannode_4_w_range4115w(0) <= atannode_4_w(20);
	wire_ccc_cordic_m_w_atannode_4_w_range4123w(0) <= atannode_4_w(21);
	wire_ccc_cordic_m_w_atannode_4_w_range4131w(0) <= atannode_4_w(22);
	wire_ccc_cordic_m_w_atannode_4_w_range4139w(0) <= atannode_4_w(23);
	wire_ccc_cordic_m_w_atannode_4_w_range4147w(0) <= atannode_4_w(24);
	wire_ccc_cordic_m_w_atannode_4_w_range4155w(0) <= atannode_4_w(25);
	wire_ccc_cordic_m_w_atannode_4_w_range4163w(0) <= atannode_4_w(26);
	wire_ccc_cordic_m_w_atannode_4_w_range4171w(0) <= atannode_4_w(27);
	wire_ccc_cordic_m_w_atannode_4_w_range4179w(0) <= atannode_4_w(28);
	wire_ccc_cordic_m_w_atannode_4_w_range4187w(0) <= atannode_4_w(29);
	wire_ccc_cordic_m_w_atannode_4_w_range3971w(0) <= atannode_4_w(2);
	wire_ccc_cordic_m_w_atannode_4_w_range4195w(0) <= atannode_4_w(30);
	wire_ccc_cordic_m_w_atannode_4_w_range4203w(0) <= atannode_4_w(31);
	wire_ccc_cordic_m_w_atannode_4_w_range4211w(0) <= atannode_4_w(32);
	wire_ccc_cordic_m_w_atannode_4_w_range4219w(0) <= atannode_4_w(33);
	wire_ccc_cordic_m_w_atannode_4_w_range3979w(0) <= atannode_4_w(3);
	wire_ccc_cordic_m_w_atannode_4_w_range3987w(0) <= atannode_4_w(4);
	wire_ccc_cordic_m_w_atannode_4_w_range3995w(0) <= atannode_4_w(5);
	wire_ccc_cordic_m_w_atannode_4_w_range4003w(0) <= atannode_4_w(6);
	wire_ccc_cordic_m_w_atannode_4_w_range4011w(0) <= atannode_4_w(7);
	wire_ccc_cordic_m_w_atannode_4_w_range4019w(0) <= atannode_4_w(8);
	wire_ccc_cordic_m_w_atannode_4_w_range4027w(0) <= atannode_4_w(9);
	wire_ccc_cordic_m_w_atannode_5_w_range4786w(0) <= atannode_5_w(0);
	wire_ccc_cordic_m_w_atannode_5_w_range4867w(0) <= atannode_5_w(10);
	wire_ccc_cordic_m_w_atannode_5_w_range4875w(0) <= atannode_5_w(11);
	wire_ccc_cordic_m_w_atannode_5_w_range4883w(0) <= atannode_5_w(12);
	wire_ccc_cordic_m_w_atannode_5_w_range4891w(0) <= atannode_5_w(13);
	wire_ccc_cordic_m_w_atannode_5_w_range4899w(0) <= atannode_5_w(14);
	wire_ccc_cordic_m_w_atannode_5_w_range4907w(0) <= atannode_5_w(15);
	wire_ccc_cordic_m_w_atannode_5_w_range4915w(0) <= atannode_5_w(16);
	wire_ccc_cordic_m_w_atannode_5_w_range4923w(0) <= atannode_5_w(17);
	wire_ccc_cordic_m_w_atannode_5_w_range4931w(0) <= atannode_5_w(18);
	wire_ccc_cordic_m_w_atannode_5_w_range4939w(0) <= atannode_5_w(19);
	wire_ccc_cordic_m_w_atannode_5_w_range4795w(0) <= atannode_5_w(1);
	wire_ccc_cordic_m_w_atannode_5_w_range4947w(0) <= atannode_5_w(20);
	wire_ccc_cordic_m_w_atannode_5_w_range4955w(0) <= atannode_5_w(21);
	wire_ccc_cordic_m_w_atannode_5_w_range4963w(0) <= atannode_5_w(22);
	wire_ccc_cordic_m_w_atannode_5_w_range4971w(0) <= atannode_5_w(23);
	wire_ccc_cordic_m_w_atannode_5_w_range4979w(0) <= atannode_5_w(24);
	wire_ccc_cordic_m_w_atannode_5_w_range4987w(0) <= atannode_5_w(25);
	wire_ccc_cordic_m_w_atannode_5_w_range4995w(0) <= atannode_5_w(26);
	wire_ccc_cordic_m_w_atannode_5_w_range5003w(0) <= atannode_5_w(27);
	wire_ccc_cordic_m_w_atannode_5_w_range5011w(0) <= atannode_5_w(28);
	wire_ccc_cordic_m_w_atannode_5_w_range5019w(0) <= atannode_5_w(29);
	wire_ccc_cordic_m_w_atannode_5_w_range4803w(0) <= atannode_5_w(2);
	wire_ccc_cordic_m_w_atannode_5_w_range5027w(0) <= atannode_5_w(30);
	wire_ccc_cordic_m_w_atannode_5_w_range5035w(0) <= atannode_5_w(31);
	wire_ccc_cordic_m_w_atannode_5_w_range5043w(0) <= atannode_5_w(32);
	wire_ccc_cordic_m_w_atannode_5_w_range5051w(0) <= atannode_5_w(33);
	wire_ccc_cordic_m_w_atannode_5_w_range4811w(0) <= atannode_5_w(3);
	wire_ccc_cordic_m_w_atannode_5_w_range4819w(0) <= atannode_5_w(4);
	wire_ccc_cordic_m_w_atannode_5_w_range4827w(0) <= atannode_5_w(5);
	wire_ccc_cordic_m_w_atannode_5_w_range4835w(0) <= atannode_5_w(6);
	wire_ccc_cordic_m_w_atannode_5_w_range4843w(0) <= atannode_5_w(7);
	wire_ccc_cordic_m_w_atannode_5_w_range4851w(0) <= atannode_5_w(8);
	wire_ccc_cordic_m_w_atannode_5_w_range4859w(0) <= atannode_5_w(9);
	wire_ccc_cordic_m_w_atannode_6_w_range5613w(0) <= atannode_6_w(0);
	wire_ccc_cordic_m_w_atannode_6_w_range5694w(0) <= atannode_6_w(10);
	wire_ccc_cordic_m_w_atannode_6_w_range5702w(0) <= atannode_6_w(11);
	wire_ccc_cordic_m_w_atannode_6_w_range5710w(0) <= atannode_6_w(12);
	wire_ccc_cordic_m_w_atannode_6_w_range5718w(0) <= atannode_6_w(13);
	wire_ccc_cordic_m_w_atannode_6_w_range5726w(0) <= atannode_6_w(14);
	wire_ccc_cordic_m_w_atannode_6_w_range5734w(0) <= atannode_6_w(15);
	wire_ccc_cordic_m_w_atannode_6_w_range5742w(0) <= atannode_6_w(16);
	wire_ccc_cordic_m_w_atannode_6_w_range5750w(0) <= atannode_6_w(17);
	wire_ccc_cordic_m_w_atannode_6_w_range5758w(0) <= atannode_6_w(18);
	wire_ccc_cordic_m_w_atannode_6_w_range5766w(0) <= atannode_6_w(19);
	wire_ccc_cordic_m_w_atannode_6_w_range5622w(0) <= atannode_6_w(1);
	wire_ccc_cordic_m_w_atannode_6_w_range5774w(0) <= atannode_6_w(20);
	wire_ccc_cordic_m_w_atannode_6_w_range5782w(0) <= atannode_6_w(21);
	wire_ccc_cordic_m_w_atannode_6_w_range5790w(0) <= atannode_6_w(22);
	wire_ccc_cordic_m_w_atannode_6_w_range5798w(0) <= atannode_6_w(23);
	wire_ccc_cordic_m_w_atannode_6_w_range5806w(0) <= atannode_6_w(24);
	wire_ccc_cordic_m_w_atannode_6_w_range5814w(0) <= atannode_6_w(25);
	wire_ccc_cordic_m_w_atannode_6_w_range5822w(0) <= atannode_6_w(26);
	wire_ccc_cordic_m_w_atannode_6_w_range5830w(0) <= atannode_6_w(27);
	wire_ccc_cordic_m_w_atannode_6_w_range5838w(0) <= atannode_6_w(28);
	wire_ccc_cordic_m_w_atannode_6_w_range5846w(0) <= atannode_6_w(29);
	wire_ccc_cordic_m_w_atannode_6_w_range5630w(0) <= atannode_6_w(2);
	wire_ccc_cordic_m_w_atannode_6_w_range5854w(0) <= atannode_6_w(30);
	wire_ccc_cordic_m_w_atannode_6_w_range5862w(0) <= atannode_6_w(31);
	wire_ccc_cordic_m_w_atannode_6_w_range5870w(0) <= atannode_6_w(32);
	wire_ccc_cordic_m_w_atannode_6_w_range5878w(0) <= atannode_6_w(33);
	wire_ccc_cordic_m_w_atannode_6_w_range5638w(0) <= atannode_6_w(3);
	wire_ccc_cordic_m_w_atannode_6_w_range5646w(0) <= atannode_6_w(4);
	wire_ccc_cordic_m_w_atannode_6_w_range5654w(0) <= atannode_6_w(5);
	wire_ccc_cordic_m_w_atannode_6_w_range5662w(0) <= atannode_6_w(6);
	wire_ccc_cordic_m_w_atannode_6_w_range5670w(0) <= atannode_6_w(7);
	wire_ccc_cordic_m_w_atannode_6_w_range5678w(0) <= atannode_6_w(8);
	wire_ccc_cordic_m_w_atannode_6_w_range5686w(0) <= atannode_6_w(9);
	wire_ccc_cordic_m_w_atannode_7_w_range6435w(0) <= atannode_7_w(0);
	wire_ccc_cordic_m_w_atannode_7_w_range6516w(0) <= atannode_7_w(10);
	wire_ccc_cordic_m_w_atannode_7_w_range6524w(0) <= atannode_7_w(11);
	wire_ccc_cordic_m_w_atannode_7_w_range6532w(0) <= atannode_7_w(12);
	wire_ccc_cordic_m_w_atannode_7_w_range6540w(0) <= atannode_7_w(13);
	wire_ccc_cordic_m_w_atannode_7_w_range6548w(0) <= atannode_7_w(14);
	wire_ccc_cordic_m_w_atannode_7_w_range6556w(0) <= atannode_7_w(15);
	wire_ccc_cordic_m_w_atannode_7_w_range6564w(0) <= atannode_7_w(16);
	wire_ccc_cordic_m_w_atannode_7_w_range6572w(0) <= atannode_7_w(17);
	wire_ccc_cordic_m_w_atannode_7_w_range6580w(0) <= atannode_7_w(18);
	wire_ccc_cordic_m_w_atannode_7_w_range6588w(0) <= atannode_7_w(19);
	wire_ccc_cordic_m_w_atannode_7_w_range6444w(0) <= atannode_7_w(1);
	wire_ccc_cordic_m_w_atannode_7_w_range6596w(0) <= atannode_7_w(20);
	wire_ccc_cordic_m_w_atannode_7_w_range6604w(0) <= atannode_7_w(21);
	wire_ccc_cordic_m_w_atannode_7_w_range6612w(0) <= atannode_7_w(22);
	wire_ccc_cordic_m_w_atannode_7_w_range6620w(0) <= atannode_7_w(23);
	wire_ccc_cordic_m_w_atannode_7_w_range6628w(0) <= atannode_7_w(24);
	wire_ccc_cordic_m_w_atannode_7_w_range6636w(0) <= atannode_7_w(25);
	wire_ccc_cordic_m_w_atannode_7_w_range6644w(0) <= atannode_7_w(26);
	wire_ccc_cordic_m_w_atannode_7_w_range6652w(0) <= atannode_7_w(27);
	wire_ccc_cordic_m_w_atannode_7_w_range6660w(0) <= atannode_7_w(28);
	wire_ccc_cordic_m_w_atannode_7_w_range6668w(0) <= atannode_7_w(29);
	wire_ccc_cordic_m_w_atannode_7_w_range6452w(0) <= atannode_7_w(2);
	wire_ccc_cordic_m_w_atannode_7_w_range6676w(0) <= atannode_7_w(30);
	wire_ccc_cordic_m_w_atannode_7_w_range6684w(0) <= atannode_7_w(31);
	wire_ccc_cordic_m_w_atannode_7_w_range6692w(0) <= atannode_7_w(32);
	wire_ccc_cordic_m_w_atannode_7_w_range6700w(0) <= atannode_7_w(33);
	wire_ccc_cordic_m_w_atannode_7_w_range6460w(0) <= atannode_7_w(3);
	wire_ccc_cordic_m_w_atannode_7_w_range6468w(0) <= atannode_7_w(4);
	wire_ccc_cordic_m_w_atannode_7_w_range6476w(0) <= atannode_7_w(5);
	wire_ccc_cordic_m_w_atannode_7_w_range6484w(0) <= atannode_7_w(6);
	wire_ccc_cordic_m_w_atannode_7_w_range6492w(0) <= atannode_7_w(7);
	wire_ccc_cordic_m_w_atannode_7_w_range6500w(0) <= atannode_7_w(8);
	wire_ccc_cordic_m_w_atannode_7_w_range6508w(0) <= atannode_7_w(9);
	wire_ccc_cordic_m_w_atannode_8_w_range7252w(0) <= atannode_8_w(0);
	wire_ccc_cordic_m_w_atannode_8_w_range7333w(0) <= atannode_8_w(10);
	wire_ccc_cordic_m_w_atannode_8_w_range7341w(0) <= atannode_8_w(11);
	wire_ccc_cordic_m_w_atannode_8_w_range7349w(0) <= atannode_8_w(12);
	wire_ccc_cordic_m_w_atannode_8_w_range7357w(0) <= atannode_8_w(13);
	wire_ccc_cordic_m_w_atannode_8_w_range7365w(0) <= atannode_8_w(14);
	wire_ccc_cordic_m_w_atannode_8_w_range7373w(0) <= atannode_8_w(15);
	wire_ccc_cordic_m_w_atannode_8_w_range7381w(0) <= atannode_8_w(16);
	wire_ccc_cordic_m_w_atannode_8_w_range7389w(0) <= atannode_8_w(17);
	wire_ccc_cordic_m_w_atannode_8_w_range7397w(0) <= atannode_8_w(18);
	wire_ccc_cordic_m_w_atannode_8_w_range7405w(0) <= atannode_8_w(19);
	wire_ccc_cordic_m_w_atannode_8_w_range7261w(0) <= atannode_8_w(1);
	wire_ccc_cordic_m_w_atannode_8_w_range7413w(0) <= atannode_8_w(20);
	wire_ccc_cordic_m_w_atannode_8_w_range7421w(0) <= atannode_8_w(21);
	wire_ccc_cordic_m_w_atannode_8_w_range7429w(0) <= atannode_8_w(22);
	wire_ccc_cordic_m_w_atannode_8_w_range7437w(0) <= atannode_8_w(23);
	wire_ccc_cordic_m_w_atannode_8_w_range7445w(0) <= atannode_8_w(24);
	wire_ccc_cordic_m_w_atannode_8_w_range7453w(0) <= atannode_8_w(25);
	wire_ccc_cordic_m_w_atannode_8_w_range7461w(0) <= atannode_8_w(26);
	wire_ccc_cordic_m_w_atannode_8_w_range7469w(0) <= atannode_8_w(27);
	wire_ccc_cordic_m_w_atannode_8_w_range7477w(0) <= atannode_8_w(28);
	wire_ccc_cordic_m_w_atannode_8_w_range7485w(0) <= atannode_8_w(29);
	wire_ccc_cordic_m_w_atannode_8_w_range7269w(0) <= atannode_8_w(2);
	wire_ccc_cordic_m_w_atannode_8_w_range7493w(0) <= atannode_8_w(30);
	wire_ccc_cordic_m_w_atannode_8_w_range7501w(0) <= atannode_8_w(31);
	wire_ccc_cordic_m_w_atannode_8_w_range7509w(0) <= atannode_8_w(32);
	wire_ccc_cordic_m_w_atannode_8_w_range7517w(0) <= atannode_8_w(33);
	wire_ccc_cordic_m_w_atannode_8_w_range7277w(0) <= atannode_8_w(3);
	wire_ccc_cordic_m_w_atannode_8_w_range7285w(0) <= atannode_8_w(4);
	wire_ccc_cordic_m_w_atannode_8_w_range7293w(0) <= atannode_8_w(5);
	wire_ccc_cordic_m_w_atannode_8_w_range7301w(0) <= atannode_8_w(6);
	wire_ccc_cordic_m_w_atannode_8_w_range7309w(0) <= atannode_8_w(7);
	wire_ccc_cordic_m_w_atannode_8_w_range7317w(0) <= atannode_8_w(8);
	wire_ccc_cordic_m_w_atannode_8_w_range7325w(0) <= atannode_8_w(9);
	wire_ccc_cordic_m_w_atannode_9_w_range8064w(0) <= atannode_9_w(0);
	wire_ccc_cordic_m_w_atannode_9_w_range8145w(0) <= atannode_9_w(10);
	wire_ccc_cordic_m_w_atannode_9_w_range8153w(0) <= atannode_9_w(11);
	wire_ccc_cordic_m_w_atannode_9_w_range8161w(0) <= atannode_9_w(12);
	wire_ccc_cordic_m_w_atannode_9_w_range8169w(0) <= atannode_9_w(13);
	wire_ccc_cordic_m_w_atannode_9_w_range8177w(0) <= atannode_9_w(14);
	wire_ccc_cordic_m_w_atannode_9_w_range8185w(0) <= atannode_9_w(15);
	wire_ccc_cordic_m_w_atannode_9_w_range8193w(0) <= atannode_9_w(16);
	wire_ccc_cordic_m_w_atannode_9_w_range8201w(0) <= atannode_9_w(17);
	wire_ccc_cordic_m_w_atannode_9_w_range8209w(0) <= atannode_9_w(18);
	wire_ccc_cordic_m_w_atannode_9_w_range8217w(0) <= atannode_9_w(19);
	wire_ccc_cordic_m_w_atannode_9_w_range8073w(0) <= atannode_9_w(1);
	wire_ccc_cordic_m_w_atannode_9_w_range8225w(0) <= atannode_9_w(20);
	wire_ccc_cordic_m_w_atannode_9_w_range8233w(0) <= atannode_9_w(21);
	wire_ccc_cordic_m_w_atannode_9_w_range8241w(0) <= atannode_9_w(22);
	wire_ccc_cordic_m_w_atannode_9_w_range8249w(0) <= atannode_9_w(23);
	wire_ccc_cordic_m_w_atannode_9_w_range8257w(0) <= atannode_9_w(24);
	wire_ccc_cordic_m_w_atannode_9_w_range8265w(0) <= atannode_9_w(25);
	wire_ccc_cordic_m_w_atannode_9_w_range8273w(0) <= atannode_9_w(26);
	wire_ccc_cordic_m_w_atannode_9_w_range8281w(0) <= atannode_9_w(27);
	wire_ccc_cordic_m_w_atannode_9_w_range8289w(0) <= atannode_9_w(28);
	wire_ccc_cordic_m_w_atannode_9_w_range8297w(0) <= atannode_9_w(29);
	wire_ccc_cordic_m_w_atannode_9_w_range8081w(0) <= atannode_9_w(2);
	wire_ccc_cordic_m_w_atannode_9_w_range8305w(0) <= atannode_9_w(30);
	wire_ccc_cordic_m_w_atannode_9_w_range8313w(0) <= atannode_9_w(31);
	wire_ccc_cordic_m_w_atannode_9_w_range8321w(0) <= atannode_9_w(32);
	wire_ccc_cordic_m_w_atannode_9_w_range8329w(0) <= atannode_9_w(33);
	wire_ccc_cordic_m_w_atannode_9_w_range8089w(0) <= atannode_9_w(3);
	wire_ccc_cordic_m_w_atannode_9_w_range8097w(0) <= atannode_9_w(4);
	wire_ccc_cordic_m_w_atannode_9_w_range8105w(0) <= atannode_9_w(5);
	wire_ccc_cordic_m_w_atannode_9_w_range8113w(0) <= atannode_9_w(6);
	wire_ccc_cordic_m_w_atannode_9_w_range8121w(0) <= atannode_9_w(7);
	wire_ccc_cordic_m_w_atannode_9_w_range8129w(0) <= atannode_9_w(8);
	wire_ccc_cordic_m_w_atannode_9_w_range8137w(0) <= atannode_9_w(9);
	wire_ccc_cordic_m_w_pre_estimate_w_range10753w(0) <= pre_estimate_w(0);
	wire_ccc_cordic_m_w_pre_estimate_w_range10794w(0) <= pre_estimate_w(10);
	wire_ccc_cordic_m_w_pre_estimate_w_range10799w(0) <= pre_estimate_w(11);
	wire_ccc_cordic_m_w_pre_estimate_w_range10804w(0) <= pre_estimate_w(12);
	wire_ccc_cordic_m_w_pre_estimate_w_range10809w(0) <= pre_estimate_w(13);
	wire_ccc_cordic_m_w_pre_estimate_w_range10814w(0) <= pre_estimate_w(14);
	wire_ccc_cordic_m_w_pre_estimate_w_range10819w(0) <= pre_estimate_w(15);
	wire_ccc_cordic_m_w_pre_estimate_w_range10824w(0) <= pre_estimate_w(16);
	wire_ccc_cordic_m_w_pre_estimate_w_range10829w(0) <= pre_estimate_w(17);
	wire_ccc_cordic_m_w_pre_estimate_w_range10834w(0) <= pre_estimate_w(18);
	wire_ccc_cordic_m_w_pre_estimate_w_range10839w(0) <= pre_estimate_w(19);
	wire_ccc_cordic_m_w_pre_estimate_w_range10760w(0) <= pre_estimate_w(1);
	wire_ccc_cordic_m_w_pre_estimate_w_range10844w(0) <= pre_estimate_w(20);
	wire_ccc_cordic_m_w_pre_estimate_w_range10849w(0) <= pre_estimate_w(21);
	wire_ccc_cordic_m_w_pre_estimate_w_range10854w(0) <= pre_estimate_w(22);
	wire_ccc_cordic_m_w_pre_estimate_w_range10859w(0) <= pre_estimate_w(23);
	wire_ccc_cordic_m_w_pre_estimate_w_range10864w(0) <= pre_estimate_w(24);
	wire_ccc_cordic_m_w_pre_estimate_w_range10869w(0) <= pre_estimate_w(25);
	wire_ccc_cordic_m_w_pre_estimate_w_range10874w(0) <= pre_estimate_w(26);
	wire_ccc_cordic_m_w_pre_estimate_w_range10879w(0) <= pre_estimate_w(27);
	wire_ccc_cordic_m_w_pre_estimate_w_range10884w(0) <= pre_estimate_w(28);
	wire_ccc_cordic_m_w_pre_estimate_w_range10889w(0) <= pre_estimate_w(29);
	wire_ccc_cordic_m_w_pre_estimate_w_range10750w(0) <= pre_estimate_w(2);
	wire_ccc_cordic_m_w_pre_estimate_w_range10894w(0) <= pre_estimate_w(30);
	wire_ccc_cordic_m_w_pre_estimate_w_range10899w(0) <= pre_estimate_w(31);
	wire_ccc_cordic_m_w_pre_estimate_w_range10904w(0) <= pre_estimate_w(32);
	wire_ccc_cordic_m_w_pre_estimate_w_range10909w(0) <= pre_estimate_w(33);
	wire_ccc_cordic_m_w_pre_estimate_w_range10758w(0) <= pre_estimate_w(3);
	wire_ccc_cordic_m_w_pre_estimate_w_range10764w(0) <= pre_estimate_w(4);
	wire_ccc_cordic_m_w_pre_estimate_w_range10769w(0) <= pre_estimate_w(5);
	wire_ccc_cordic_m_w_pre_estimate_w_range10774w(0) <= pre_estimate_w(6);
	wire_ccc_cordic_m_w_pre_estimate_w_range10779w(0) <= pre_estimate_w(7);
	wire_ccc_cordic_m_w_pre_estimate_w_range10784w(0) <= pre_estimate_w(8);
	wire_ccc_cordic_m_w_pre_estimate_w_range10789w(0) <= pre_estimate_w(9);
	wire_ccc_cordic_m_w_radians_range410w(0) <= radians(0);
	wire_ccc_cordic_m_w_radians_range458w(0) <= radians(10);
	wire_ccc_cordic_m_w_radians_range463w(0) <= radians(11);
	wire_ccc_cordic_m_w_radians_range468w(0) <= radians(12);
	wire_ccc_cordic_m_w_radians_range473w(0) <= radians(13);
	wire_ccc_cordic_m_w_radians_range478w(0) <= radians(14);
	wire_ccc_cordic_m_w_radians_range483w(0) <= radians(15);
	wire_ccc_cordic_m_w_radians_range488w(0) <= radians(16);
	wire_ccc_cordic_m_w_radians_range493w(0) <= radians(17);
	wire_ccc_cordic_m_w_radians_range498w(0) <= radians(18);
	wire_ccc_cordic_m_w_radians_range503w(0) <= radians(19);
	wire_ccc_cordic_m_w_radians_range415w(0) <= radians(1);
	wire_ccc_cordic_m_w_radians_range508w(0) <= radians(20);
	wire_ccc_cordic_m_w_radians_range513w(0) <= radians(21);
	wire_ccc_cordic_m_w_radians_range518w(0) <= radians(22);
	wire_ccc_cordic_m_w_radians_range523w(0) <= radians(23);
	wire_ccc_cordic_m_w_radians_range528w(0) <= radians(24);
	wire_ccc_cordic_m_w_radians_range533w(0) <= radians(25);
	wire_ccc_cordic_m_w_radians_range538w(0) <= radians(26);
	wire_ccc_cordic_m_w_radians_range543w(0) <= radians(27);
	wire_ccc_cordic_m_w_radians_range548w(0) <= radians(28);
	wire_ccc_cordic_m_w_radians_range553w(0) <= radians(29);
	wire_ccc_cordic_m_w_radians_range418w(0) <= radians(2);
	wire_ccc_cordic_m_w_radians_range558w(0) <= radians(30);
	wire_ccc_cordic_m_w_radians_range563w(0) <= radians(31);
	wire_ccc_cordic_m_w_radians_range568w(0) <= radians(32);
	wire_ccc_cordic_m_w_radians_range573w(0) <= radians(33);
	wire_ccc_cordic_m_w_radians_range423w(0) <= radians(3);
	wire_ccc_cordic_m_w_radians_range428w(0) <= radians(4);
	wire_ccc_cordic_m_w_radians_range433w(0) <= radians(5);
	wire_ccc_cordic_m_w_radians_range438w(0) <= radians(6);
	wire_ccc_cordic_m_w_radians_range443w(0) <= radians(7);
	wire_ccc_cordic_m_w_radians_range448w(0) <= radians(8);
	wire_ccc_cordic_m_w_radians_range453w(0) <= radians(9);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7786w(0) <= x_prenode_10_w(0);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7868w(0) <= x_prenode_10_w(10);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7876w(0) <= x_prenode_10_w(11);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7884w(0) <= x_prenode_10_w(12);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7892w(0) <= x_prenode_10_w(13);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7900w(0) <= x_prenode_10_w(14);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7908w(0) <= x_prenode_10_w(15);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7916w(0) <= x_prenode_10_w(16);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7924w(0) <= x_prenode_10_w(17);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7932w(0) <= x_prenode_10_w(18);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7940w(0) <= x_prenode_10_w(19);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7796w(0) <= x_prenode_10_w(1);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7948w(0) <= x_prenode_10_w(20);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7956w(0) <= x_prenode_10_w(21);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7964w(0) <= x_prenode_10_w(22);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7972w(0) <= x_prenode_10_w(23);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7980w(0) <= x_prenode_10_w(24);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7988w(0) <= x_prenode_10_w(25);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7996w(0) <= x_prenode_10_w(26);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8004w(0) <= x_prenode_10_w(27);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8012w(0) <= x_prenode_10_w(28);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8020w(0) <= x_prenode_10_w(29);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7804w(0) <= x_prenode_10_w(2);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8028w(0) <= x_prenode_10_w(30);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8036w(0) <= x_prenode_10_w(31);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8044w(0) <= x_prenode_10_w(32);
	wire_ccc_cordic_m_w_x_prenode_10_w_range8052w(0) <= x_prenode_10_w(33);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7812w(0) <= x_prenode_10_w(3);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7820w(0) <= x_prenode_10_w(4);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7828w(0) <= x_prenode_10_w(5);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7836w(0) <= x_prenode_10_w(6);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7844w(0) <= x_prenode_10_w(7);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7852w(0) <= x_prenode_10_w(8);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7860w(0) <= x_prenode_10_w(9);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8593w(0) <= x_prenode_11_w(0);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8675w(0) <= x_prenode_11_w(10);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8683w(0) <= x_prenode_11_w(11);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8691w(0) <= x_prenode_11_w(12);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8699w(0) <= x_prenode_11_w(13);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8707w(0) <= x_prenode_11_w(14);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8715w(0) <= x_prenode_11_w(15);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8723w(0) <= x_prenode_11_w(16);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8731w(0) <= x_prenode_11_w(17);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8739w(0) <= x_prenode_11_w(18);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8747w(0) <= x_prenode_11_w(19);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8603w(0) <= x_prenode_11_w(1);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8755w(0) <= x_prenode_11_w(20);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8763w(0) <= x_prenode_11_w(21);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8771w(0) <= x_prenode_11_w(22);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8779w(0) <= x_prenode_11_w(23);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8787w(0) <= x_prenode_11_w(24);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8795w(0) <= x_prenode_11_w(25);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8803w(0) <= x_prenode_11_w(26);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8811w(0) <= x_prenode_11_w(27);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8819w(0) <= x_prenode_11_w(28);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8827w(0) <= x_prenode_11_w(29);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8611w(0) <= x_prenode_11_w(2);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8835w(0) <= x_prenode_11_w(30);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8843w(0) <= x_prenode_11_w(31);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8851w(0) <= x_prenode_11_w(32);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8859w(0) <= x_prenode_11_w(33);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8619w(0) <= x_prenode_11_w(3);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8627w(0) <= x_prenode_11_w(4);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8635w(0) <= x_prenode_11_w(5);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8643w(0) <= x_prenode_11_w(6);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8651w(0) <= x_prenode_11_w(7);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8659w(0) <= x_prenode_11_w(8);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8667w(0) <= x_prenode_11_w(9);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9395w(0) <= x_prenode_12_w(0);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9477w(0) <= x_prenode_12_w(10);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9485w(0) <= x_prenode_12_w(11);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9493w(0) <= x_prenode_12_w(12);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9501w(0) <= x_prenode_12_w(13);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9509w(0) <= x_prenode_12_w(14);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9517w(0) <= x_prenode_12_w(15);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9525w(0) <= x_prenode_12_w(16);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9533w(0) <= x_prenode_12_w(17);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9541w(0) <= x_prenode_12_w(18);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9549w(0) <= x_prenode_12_w(19);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9405w(0) <= x_prenode_12_w(1);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9557w(0) <= x_prenode_12_w(20);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9565w(0) <= x_prenode_12_w(21);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9573w(0) <= x_prenode_12_w(22);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9581w(0) <= x_prenode_12_w(23);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9589w(0) <= x_prenode_12_w(24);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9597w(0) <= x_prenode_12_w(25);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9605w(0) <= x_prenode_12_w(26);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9613w(0) <= x_prenode_12_w(27);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9621w(0) <= x_prenode_12_w(28);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9629w(0) <= x_prenode_12_w(29);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9413w(0) <= x_prenode_12_w(2);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9637w(0) <= x_prenode_12_w(30);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9645w(0) <= x_prenode_12_w(31);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9653w(0) <= x_prenode_12_w(32);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9661w(0) <= x_prenode_12_w(33);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9421w(0) <= x_prenode_12_w(3);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9429w(0) <= x_prenode_12_w(4);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9437w(0) <= x_prenode_12_w(5);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9445w(0) <= x_prenode_12_w(6);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9453w(0) <= x_prenode_12_w(7);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9461w(0) <= x_prenode_12_w(8);
	wire_ccc_cordic_m_w_x_prenode_12_w_range9469w(0) <= x_prenode_12_w(9);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10192w(0) <= x_prenode_13_w(0);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10274w(0) <= x_prenode_13_w(10);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10282w(0) <= x_prenode_13_w(11);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10290w(0) <= x_prenode_13_w(12);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10298w(0) <= x_prenode_13_w(13);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10306w(0) <= x_prenode_13_w(14);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10314w(0) <= x_prenode_13_w(15);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10322w(0) <= x_prenode_13_w(16);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10330w(0) <= x_prenode_13_w(17);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10338w(0) <= x_prenode_13_w(18);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10346w(0) <= x_prenode_13_w(19);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10202w(0) <= x_prenode_13_w(1);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10354w(0) <= x_prenode_13_w(20);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10362w(0) <= x_prenode_13_w(21);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10370w(0) <= x_prenode_13_w(22);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10378w(0) <= x_prenode_13_w(23);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10386w(0) <= x_prenode_13_w(24);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10394w(0) <= x_prenode_13_w(25);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10402w(0) <= x_prenode_13_w(26);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10410w(0) <= x_prenode_13_w(27);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10418w(0) <= x_prenode_13_w(28);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10426w(0) <= x_prenode_13_w(29);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10210w(0) <= x_prenode_13_w(2);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10434w(0) <= x_prenode_13_w(30);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10442w(0) <= x_prenode_13_w(31);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10450w(0) <= x_prenode_13_w(32);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10458w(0) <= x_prenode_13_w(33);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10218w(0) <= x_prenode_13_w(3);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10226w(0) <= x_prenode_13_w(4);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10234w(0) <= x_prenode_13_w(5);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10242w(0) <= x_prenode_13_w(6);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10250w(0) <= x_prenode_13_w(7);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10258w(0) <= x_prenode_13_w(8);
	wire_ccc_cordic_m_w_x_prenode_13_w_range10266w(0) <= x_prenode_13_w(9);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1150w(0) <= x_prenode_2_w(0);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1232w(0) <= x_prenode_2_w(10);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1240w(0) <= x_prenode_2_w(11);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1248w(0) <= x_prenode_2_w(12);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1256w(0) <= x_prenode_2_w(13);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1264w(0) <= x_prenode_2_w(14);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1272w(0) <= x_prenode_2_w(15);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1280w(0) <= x_prenode_2_w(16);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1288w(0) <= x_prenode_2_w(17);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1296w(0) <= x_prenode_2_w(18);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1304w(0) <= x_prenode_2_w(19);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1160w(0) <= x_prenode_2_w(1);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1312w(0) <= x_prenode_2_w(20);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1320w(0) <= x_prenode_2_w(21);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1328w(0) <= x_prenode_2_w(22);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1336w(0) <= x_prenode_2_w(23);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1344w(0) <= x_prenode_2_w(24);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1352w(0) <= x_prenode_2_w(25);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1360w(0) <= x_prenode_2_w(26);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1368w(0) <= x_prenode_2_w(27);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1376w(0) <= x_prenode_2_w(28);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1384w(0) <= x_prenode_2_w(29);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1168w(0) <= x_prenode_2_w(2);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1392w(0) <= x_prenode_2_w(30);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1400w(0) <= x_prenode_2_w(31);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1408w(0) <= x_prenode_2_w(32);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1416w(0) <= x_prenode_2_w(33);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1176w(0) <= x_prenode_2_w(3);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1184w(0) <= x_prenode_2_w(4);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1192w(0) <= x_prenode_2_w(5);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1200w(0) <= x_prenode_2_w(6);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1208w(0) <= x_prenode_2_w(7);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1216w(0) <= x_prenode_2_w(8);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1224w(0) <= x_prenode_2_w(9);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1997w(0) <= x_prenode_3_w(0);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2079w(0) <= x_prenode_3_w(10);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2087w(0) <= x_prenode_3_w(11);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2095w(0) <= x_prenode_3_w(12);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2103w(0) <= x_prenode_3_w(13);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2111w(0) <= x_prenode_3_w(14);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2119w(0) <= x_prenode_3_w(15);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2127w(0) <= x_prenode_3_w(16);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2135w(0) <= x_prenode_3_w(17);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2143w(0) <= x_prenode_3_w(18);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2151w(0) <= x_prenode_3_w(19);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2007w(0) <= x_prenode_3_w(1);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2159w(0) <= x_prenode_3_w(20);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2167w(0) <= x_prenode_3_w(21);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2175w(0) <= x_prenode_3_w(22);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2183w(0) <= x_prenode_3_w(23);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2191w(0) <= x_prenode_3_w(24);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2199w(0) <= x_prenode_3_w(25);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2207w(0) <= x_prenode_3_w(26);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2215w(0) <= x_prenode_3_w(27);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2223w(0) <= x_prenode_3_w(28);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2231w(0) <= x_prenode_3_w(29);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2015w(0) <= x_prenode_3_w(2);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2239w(0) <= x_prenode_3_w(30);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2247w(0) <= x_prenode_3_w(31);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2255w(0) <= x_prenode_3_w(32);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2263w(0) <= x_prenode_3_w(33);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2023w(0) <= x_prenode_3_w(3);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2031w(0) <= x_prenode_3_w(4);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2039w(0) <= x_prenode_3_w(5);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2047w(0) <= x_prenode_3_w(6);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2055w(0) <= x_prenode_3_w(7);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2063w(0) <= x_prenode_3_w(8);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2071w(0) <= x_prenode_3_w(9);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2839w(0) <= x_prenode_4_w(0);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2921w(0) <= x_prenode_4_w(10);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2929w(0) <= x_prenode_4_w(11);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2937w(0) <= x_prenode_4_w(12);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2945w(0) <= x_prenode_4_w(13);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2953w(0) <= x_prenode_4_w(14);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2961w(0) <= x_prenode_4_w(15);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2969w(0) <= x_prenode_4_w(16);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2977w(0) <= x_prenode_4_w(17);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2985w(0) <= x_prenode_4_w(18);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2993w(0) <= x_prenode_4_w(19);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2849w(0) <= x_prenode_4_w(1);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3001w(0) <= x_prenode_4_w(20);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3009w(0) <= x_prenode_4_w(21);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3017w(0) <= x_prenode_4_w(22);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3025w(0) <= x_prenode_4_w(23);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3033w(0) <= x_prenode_4_w(24);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3041w(0) <= x_prenode_4_w(25);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3049w(0) <= x_prenode_4_w(26);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3057w(0) <= x_prenode_4_w(27);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3065w(0) <= x_prenode_4_w(28);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3073w(0) <= x_prenode_4_w(29);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2857w(0) <= x_prenode_4_w(2);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3081w(0) <= x_prenode_4_w(30);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3089w(0) <= x_prenode_4_w(31);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3097w(0) <= x_prenode_4_w(32);
	wire_ccc_cordic_m_w_x_prenode_4_w_range3105w(0) <= x_prenode_4_w(33);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2865w(0) <= x_prenode_4_w(3);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2873w(0) <= x_prenode_4_w(4);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2881w(0) <= x_prenode_4_w(5);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2889w(0) <= x_prenode_4_w(6);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2897w(0) <= x_prenode_4_w(7);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2905w(0) <= x_prenode_4_w(8);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2913w(0) <= x_prenode_4_w(9);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3676w(0) <= x_prenode_5_w(0);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3758w(0) <= x_prenode_5_w(10);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3766w(0) <= x_prenode_5_w(11);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3774w(0) <= x_prenode_5_w(12);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3782w(0) <= x_prenode_5_w(13);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3790w(0) <= x_prenode_5_w(14);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3798w(0) <= x_prenode_5_w(15);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3806w(0) <= x_prenode_5_w(16);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3814w(0) <= x_prenode_5_w(17);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3822w(0) <= x_prenode_5_w(18);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3830w(0) <= x_prenode_5_w(19);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3686w(0) <= x_prenode_5_w(1);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3838w(0) <= x_prenode_5_w(20);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3846w(0) <= x_prenode_5_w(21);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3854w(0) <= x_prenode_5_w(22);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3862w(0) <= x_prenode_5_w(23);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3870w(0) <= x_prenode_5_w(24);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3878w(0) <= x_prenode_5_w(25);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3886w(0) <= x_prenode_5_w(26);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3894w(0) <= x_prenode_5_w(27);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3902w(0) <= x_prenode_5_w(28);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3910w(0) <= x_prenode_5_w(29);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3694w(0) <= x_prenode_5_w(2);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3918w(0) <= x_prenode_5_w(30);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3926w(0) <= x_prenode_5_w(31);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3934w(0) <= x_prenode_5_w(32);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3942w(0) <= x_prenode_5_w(33);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3702w(0) <= x_prenode_5_w(3);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3710w(0) <= x_prenode_5_w(4);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3718w(0) <= x_prenode_5_w(5);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3726w(0) <= x_prenode_5_w(6);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3734w(0) <= x_prenode_5_w(7);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3742w(0) <= x_prenode_5_w(8);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3750w(0) <= x_prenode_5_w(9);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4508w(0) <= x_prenode_6_w(0);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4590w(0) <= x_prenode_6_w(10);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4598w(0) <= x_prenode_6_w(11);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4606w(0) <= x_prenode_6_w(12);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4614w(0) <= x_prenode_6_w(13);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4622w(0) <= x_prenode_6_w(14);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4630w(0) <= x_prenode_6_w(15);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4638w(0) <= x_prenode_6_w(16);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4646w(0) <= x_prenode_6_w(17);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4654w(0) <= x_prenode_6_w(18);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4662w(0) <= x_prenode_6_w(19);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4518w(0) <= x_prenode_6_w(1);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4670w(0) <= x_prenode_6_w(20);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4678w(0) <= x_prenode_6_w(21);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4686w(0) <= x_prenode_6_w(22);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4694w(0) <= x_prenode_6_w(23);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4702w(0) <= x_prenode_6_w(24);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4710w(0) <= x_prenode_6_w(25);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4718w(0) <= x_prenode_6_w(26);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4726w(0) <= x_prenode_6_w(27);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4734w(0) <= x_prenode_6_w(28);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4742w(0) <= x_prenode_6_w(29);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4526w(0) <= x_prenode_6_w(2);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4750w(0) <= x_prenode_6_w(30);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4758w(0) <= x_prenode_6_w(31);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4766w(0) <= x_prenode_6_w(32);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4774w(0) <= x_prenode_6_w(33);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4534w(0) <= x_prenode_6_w(3);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4542w(0) <= x_prenode_6_w(4);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4550w(0) <= x_prenode_6_w(5);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4558w(0) <= x_prenode_6_w(6);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4566w(0) <= x_prenode_6_w(7);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4574w(0) <= x_prenode_6_w(8);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4582w(0) <= x_prenode_6_w(9);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5335w(0) <= x_prenode_7_w(0);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5417w(0) <= x_prenode_7_w(10);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5425w(0) <= x_prenode_7_w(11);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5433w(0) <= x_prenode_7_w(12);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5441w(0) <= x_prenode_7_w(13);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5449w(0) <= x_prenode_7_w(14);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5457w(0) <= x_prenode_7_w(15);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5465w(0) <= x_prenode_7_w(16);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5473w(0) <= x_prenode_7_w(17);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5481w(0) <= x_prenode_7_w(18);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5489w(0) <= x_prenode_7_w(19);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5345w(0) <= x_prenode_7_w(1);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5497w(0) <= x_prenode_7_w(20);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5505w(0) <= x_prenode_7_w(21);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5513w(0) <= x_prenode_7_w(22);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5521w(0) <= x_prenode_7_w(23);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5529w(0) <= x_prenode_7_w(24);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5537w(0) <= x_prenode_7_w(25);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5545w(0) <= x_prenode_7_w(26);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5553w(0) <= x_prenode_7_w(27);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5561w(0) <= x_prenode_7_w(28);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5569w(0) <= x_prenode_7_w(29);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5353w(0) <= x_prenode_7_w(2);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5577w(0) <= x_prenode_7_w(30);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5585w(0) <= x_prenode_7_w(31);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5593w(0) <= x_prenode_7_w(32);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5601w(0) <= x_prenode_7_w(33);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5361w(0) <= x_prenode_7_w(3);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5369w(0) <= x_prenode_7_w(4);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5377w(0) <= x_prenode_7_w(5);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5385w(0) <= x_prenode_7_w(6);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5393w(0) <= x_prenode_7_w(7);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5401w(0) <= x_prenode_7_w(8);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5409w(0) <= x_prenode_7_w(9);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6157w(0) <= x_prenode_8_w(0);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6239w(0) <= x_prenode_8_w(10);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6247w(0) <= x_prenode_8_w(11);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6255w(0) <= x_prenode_8_w(12);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6263w(0) <= x_prenode_8_w(13);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6271w(0) <= x_prenode_8_w(14);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6279w(0) <= x_prenode_8_w(15);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6287w(0) <= x_prenode_8_w(16);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6295w(0) <= x_prenode_8_w(17);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6303w(0) <= x_prenode_8_w(18);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6311w(0) <= x_prenode_8_w(19);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6167w(0) <= x_prenode_8_w(1);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6319w(0) <= x_prenode_8_w(20);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6327w(0) <= x_prenode_8_w(21);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6335w(0) <= x_prenode_8_w(22);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6343w(0) <= x_prenode_8_w(23);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6351w(0) <= x_prenode_8_w(24);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6359w(0) <= x_prenode_8_w(25);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6367w(0) <= x_prenode_8_w(26);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6375w(0) <= x_prenode_8_w(27);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6383w(0) <= x_prenode_8_w(28);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6391w(0) <= x_prenode_8_w(29);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6175w(0) <= x_prenode_8_w(2);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6399w(0) <= x_prenode_8_w(30);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6407w(0) <= x_prenode_8_w(31);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6415w(0) <= x_prenode_8_w(32);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6423w(0) <= x_prenode_8_w(33);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6183w(0) <= x_prenode_8_w(3);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6191w(0) <= x_prenode_8_w(4);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6199w(0) <= x_prenode_8_w(5);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6207w(0) <= x_prenode_8_w(6);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6215w(0) <= x_prenode_8_w(7);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6223w(0) <= x_prenode_8_w(8);
	wire_ccc_cordic_m_w_x_prenode_8_w_range6231w(0) <= x_prenode_8_w(9);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6974w(0) <= x_prenode_9_w(0);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7056w(0) <= x_prenode_9_w(10);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7064w(0) <= x_prenode_9_w(11);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7072w(0) <= x_prenode_9_w(12);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7080w(0) <= x_prenode_9_w(13);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7088w(0) <= x_prenode_9_w(14);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7096w(0) <= x_prenode_9_w(15);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7104w(0) <= x_prenode_9_w(16);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7112w(0) <= x_prenode_9_w(17);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7120w(0) <= x_prenode_9_w(18);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7128w(0) <= x_prenode_9_w(19);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6984w(0) <= x_prenode_9_w(1);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7136w(0) <= x_prenode_9_w(20);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7144w(0) <= x_prenode_9_w(21);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7152w(0) <= x_prenode_9_w(22);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7160w(0) <= x_prenode_9_w(23);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7168w(0) <= x_prenode_9_w(24);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7176w(0) <= x_prenode_9_w(25);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7184w(0) <= x_prenode_9_w(26);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7192w(0) <= x_prenode_9_w(27);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7200w(0) <= x_prenode_9_w(28);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7208w(0) <= x_prenode_9_w(29);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6992w(0) <= x_prenode_9_w(2);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7216w(0) <= x_prenode_9_w(30);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7224w(0) <= x_prenode_9_w(31);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7232w(0) <= x_prenode_9_w(32);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7240w(0) <= x_prenode_9_w(33);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7000w(0) <= x_prenode_9_w(3);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7008w(0) <= x_prenode_9_w(4);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7016w(0) <= x_prenode_9_w(5);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7024w(0) <= x_prenode_9_w(6);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7032w(0) <= x_prenode_9_w(7);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7040w(0) <= x_prenode_9_w(8);
	wire_ccc_cordic_m_w_x_prenode_9_w_range7048w(0) <= x_prenode_9_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7570w(0) <= x_prenodeone_10_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7629w(0) <= x_prenodeone_10_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7635w(0) <= x_prenodeone_10_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7641w(0) <= x_prenodeone_10_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7647w(0) <= x_prenodeone_10_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7653w(0) <= x_prenodeone_10_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7659w(0) <= x_prenodeone_10_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7665w(0) <= x_prenodeone_10_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7671w(0) <= x_prenodeone_10_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7677w(0) <= x_prenodeone_10_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7683w(0) <= x_prenodeone_10_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7575w(0) <= x_prenodeone_10_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7689w(0) <= x_prenodeone_10_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7695w(0) <= x_prenodeone_10_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7701w(0) <= x_prenodeone_10_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7707w(0) <= x_prenodeone_10_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7711w(0) <= x_prenodeone_10_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7523w(0) <= x_prenodeone_10_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7528w(0) <= x_prenodeone_10_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7530w(0) <= x_prenodeone_10_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7532w(0) <= x_prenodeone_10_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7534w(0) <= x_prenodeone_10_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7581w(0) <= x_prenodeone_10_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7536w(0) <= x_prenodeone_10_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7538w(0) <= x_prenodeone_10_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7540w(0) <= x_prenodeone_10_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7542w(0) <= x_prenodeone_10_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7587w(0) <= x_prenodeone_10_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7593w(0) <= x_prenodeone_10_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7599w(0) <= x_prenodeone_10_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7605w(0) <= x_prenodeone_10_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7611w(0) <= x_prenodeone_10_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7617w(0) <= x_prenodeone_10_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7623w(0) <= x_prenodeone_10_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8386w(0) <= x_prenodeone_11_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8445w(0) <= x_prenodeone_11_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8451w(0) <= x_prenodeone_11_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8457w(0) <= x_prenodeone_11_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8463w(0) <= x_prenodeone_11_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8469w(0) <= x_prenodeone_11_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8475w(0) <= x_prenodeone_11_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8481w(0) <= x_prenodeone_11_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8487w(0) <= x_prenodeone_11_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8493w(0) <= x_prenodeone_11_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8499w(0) <= x_prenodeone_11_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8391w(0) <= x_prenodeone_11_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8505w(0) <= x_prenodeone_11_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8511w(0) <= x_prenodeone_11_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8517w(0) <= x_prenodeone_11_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8521w(0) <= x_prenodeone_11_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8335w(0) <= x_prenodeone_11_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8340w(0) <= x_prenodeone_11_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8342w(0) <= x_prenodeone_11_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8344w(0) <= x_prenodeone_11_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8346w(0) <= x_prenodeone_11_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8348w(0) <= x_prenodeone_11_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8397w(0) <= x_prenodeone_11_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8350w(0) <= x_prenodeone_11_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8352w(0) <= x_prenodeone_11_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8354w(0) <= x_prenodeone_11_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8356w(0) <= x_prenodeone_11_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8403w(0) <= x_prenodeone_11_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8409w(0) <= x_prenodeone_11_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8415w(0) <= x_prenodeone_11_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8421w(0) <= x_prenodeone_11_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8427w(0) <= x_prenodeone_11_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8433w(0) <= x_prenodeone_11_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range8439w(0) <= x_prenodeone_11_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9197w(0) <= x_prenodeone_12_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9256w(0) <= x_prenodeone_12_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9262w(0) <= x_prenodeone_12_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9268w(0) <= x_prenodeone_12_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9274w(0) <= x_prenodeone_12_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9280w(0) <= x_prenodeone_12_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9286w(0) <= x_prenodeone_12_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9292w(0) <= x_prenodeone_12_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9298w(0) <= x_prenodeone_12_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9304w(0) <= x_prenodeone_12_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9310w(0) <= x_prenodeone_12_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9202w(0) <= x_prenodeone_12_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9316w(0) <= x_prenodeone_12_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9322w(0) <= x_prenodeone_12_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9326w(0) <= x_prenodeone_12_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9142w(0) <= x_prenodeone_12_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9147w(0) <= x_prenodeone_12_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9149w(0) <= x_prenodeone_12_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9151w(0) <= x_prenodeone_12_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9153w(0) <= x_prenodeone_12_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9155w(0) <= x_prenodeone_12_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9157w(0) <= x_prenodeone_12_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9208w(0) <= x_prenodeone_12_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9159w(0) <= x_prenodeone_12_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9161w(0) <= x_prenodeone_12_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9163w(0) <= x_prenodeone_12_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9165w(0) <= x_prenodeone_12_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9214w(0) <= x_prenodeone_12_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9220w(0) <= x_prenodeone_12_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9226w(0) <= x_prenodeone_12_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9232w(0) <= x_prenodeone_12_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9238w(0) <= x_prenodeone_12_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9244w(0) <= x_prenodeone_12_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range9250w(0) <= x_prenodeone_12_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10003w(0) <= x_prenodeone_13_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10062w(0) <= x_prenodeone_13_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10068w(0) <= x_prenodeone_13_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10074w(0) <= x_prenodeone_13_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10080w(0) <= x_prenodeone_13_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10086w(0) <= x_prenodeone_13_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10092w(0) <= x_prenodeone_13_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10098w(0) <= x_prenodeone_13_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10104w(0) <= x_prenodeone_13_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10110w(0) <= x_prenodeone_13_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10116w(0) <= x_prenodeone_13_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10008w(0) <= x_prenodeone_13_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10122w(0) <= x_prenodeone_13_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10126w(0) <= x_prenodeone_13_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9944w(0) <= x_prenodeone_13_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9949w(0) <= x_prenodeone_13_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9951w(0) <= x_prenodeone_13_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9953w(0) <= x_prenodeone_13_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9955w(0) <= x_prenodeone_13_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9957w(0) <= x_prenodeone_13_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9959w(0) <= x_prenodeone_13_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9961w(0) <= x_prenodeone_13_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10014w(0) <= x_prenodeone_13_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9963w(0) <= x_prenodeone_13_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9965w(0) <= x_prenodeone_13_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9967w(0) <= x_prenodeone_13_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9969w(0) <= x_prenodeone_13_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10020w(0) <= x_prenodeone_13_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10026w(0) <= x_prenodeone_13_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10032w(0) <= x_prenodeone_13_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10038w(0) <= x_prenodeone_13_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10044w(0) <= x_prenodeone_13_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10050w(0) <= x_prenodeone_13_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range10056w(0) <= x_prenodeone_13_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range862w(0) <= x_prenodeone_2_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range921w(0) <= x_prenodeone_2_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range927w(0) <= x_prenodeone_2_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range933w(0) <= x_prenodeone_2_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range939w(0) <= x_prenodeone_2_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range945w(0) <= x_prenodeone_2_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range951w(0) <= x_prenodeone_2_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range957w(0) <= x_prenodeone_2_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range963w(0) <= x_prenodeone_2_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range969w(0) <= x_prenodeone_2_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range975w(0) <= x_prenodeone_2_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range867w(0) <= x_prenodeone_2_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range981w(0) <= x_prenodeone_2_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range987w(0) <= x_prenodeone_2_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range993w(0) <= x_prenodeone_2_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range999w(0) <= x_prenodeone_2_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1005w(0) <= x_prenodeone_2_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1011w(0) <= x_prenodeone_2_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1017w(0) <= x_prenodeone_2_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1023w(0) <= x_prenodeone_2_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1029w(0) <= x_prenodeone_2_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1035w(0) <= x_prenodeone_2_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range873w(0) <= x_prenodeone_2_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1041w(0) <= x_prenodeone_2_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1047w(0) <= x_prenodeone_2_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range1051w(0) <= x_prenodeone_2_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range847w(0) <= x_prenodeone_2_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range879w(0) <= x_prenodeone_2_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range885w(0) <= x_prenodeone_2_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range891w(0) <= x_prenodeone_2_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range897w(0) <= x_prenodeone_2_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range903w(0) <= x_prenodeone_2_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range909w(0) <= x_prenodeone_2_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range915w(0) <= x_prenodeone_2_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1718w(0) <= x_prenodeone_3_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1777w(0) <= x_prenodeone_3_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1783w(0) <= x_prenodeone_3_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1789w(0) <= x_prenodeone_3_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1795w(0) <= x_prenodeone_3_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1801w(0) <= x_prenodeone_3_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1807w(0) <= x_prenodeone_3_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1813w(0) <= x_prenodeone_3_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1819w(0) <= x_prenodeone_3_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1825w(0) <= x_prenodeone_3_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1831w(0) <= x_prenodeone_3_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1723w(0) <= x_prenodeone_3_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1837w(0) <= x_prenodeone_3_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1843w(0) <= x_prenodeone_3_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1849w(0) <= x_prenodeone_3_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1855w(0) <= x_prenodeone_3_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1861w(0) <= x_prenodeone_3_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1867w(0) <= x_prenodeone_3_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1873w(0) <= x_prenodeone_3_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1879w(0) <= x_prenodeone_3_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1885w(0) <= x_prenodeone_3_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1891w(0) <= x_prenodeone_3_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1729w(0) <= x_prenodeone_3_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1897w(0) <= x_prenodeone_3_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1901w(0) <= x_prenodeone_3_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1699w(0) <= x_prenodeone_3_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1704w(0) <= x_prenodeone_3_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1735w(0) <= x_prenodeone_3_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1741w(0) <= x_prenodeone_3_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1747w(0) <= x_prenodeone_3_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1753w(0) <= x_prenodeone_3_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1759w(0) <= x_prenodeone_3_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1765w(0) <= x_prenodeone_3_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1771w(0) <= x_prenodeone_3_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2569w(0) <= x_prenodeone_4_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2628w(0) <= x_prenodeone_4_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2634w(0) <= x_prenodeone_4_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2640w(0) <= x_prenodeone_4_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2646w(0) <= x_prenodeone_4_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2652w(0) <= x_prenodeone_4_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2658w(0) <= x_prenodeone_4_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2664w(0) <= x_prenodeone_4_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2670w(0) <= x_prenodeone_4_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2676w(0) <= x_prenodeone_4_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2682w(0) <= x_prenodeone_4_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2574w(0) <= x_prenodeone_4_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2688w(0) <= x_prenodeone_4_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2694w(0) <= x_prenodeone_4_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2700w(0) <= x_prenodeone_4_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2706w(0) <= x_prenodeone_4_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2712w(0) <= x_prenodeone_4_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2718w(0) <= x_prenodeone_4_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2724w(0) <= x_prenodeone_4_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2730w(0) <= x_prenodeone_4_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2736w(0) <= x_prenodeone_4_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2742w(0) <= x_prenodeone_4_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2580w(0) <= x_prenodeone_4_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2746w(0) <= x_prenodeone_4_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2546w(0) <= x_prenodeone_4_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2551w(0) <= x_prenodeone_4_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2553w(0) <= x_prenodeone_4_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2586w(0) <= x_prenodeone_4_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2592w(0) <= x_prenodeone_4_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2598w(0) <= x_prenodeone_4_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2604w(0) <= x_prenodeone_4_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2610w(0) <= x_prenodeone_4_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2616w(0) <= x_prenodeone_4_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2622w(0) <= x_prenodeone_4_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3415w(0) <= x_prenodeone_5_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3474w(0) <= x_prenodeone_5_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3480w(0) <= x_prenodeone_5_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3486w(0) <= x_prenodeone_5_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3492w(0) <= x_prenodeone_5_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3498w(0) <= x_prenodeone_5_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3504w(0) <= x_prenodeone_5_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3510w(0) <= x_prenodeone_5_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3516w(0) <= x_prenodeone_5_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3522w(0) <= x_prenodeone_5_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3528w(0) <= x_prenodeone_5_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3420w(0) <= x_prenodeone_5_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3534w(0) <= x_prenodeone_5_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3540w(0) <= x_prenodeone_5_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3546w(0) <= x_prenodeone_5_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3552w(0) <= x_prenodeone_5_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3558w(0) <= x_prenodeone_5_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3564w(0) <= x_prenodeone_5_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3570w(0) <= x_prenodeone_5_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3576w(0) <= x_prenodeone_5_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3582w(0) <= x_prenodeone_5_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3586w(0) <= x_prenodeone_5_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3426w(0) <= x_prenodeone_5_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3388w(0) <= x_prenodeone_5_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3393w(0) <= x_prenodeone_5_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3395w(0) <= x_prenodeone_5_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3397w(0) <= x_prenodeone_5_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3432w(0) <= x_prenodeone_5_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3438w(0) <= x_prenodeone_5_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3444w(0) <= x_prenodeone_5_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3450w(0) <= x_prenodeone_5_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3456w(0) <= x_prenodeone_5_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3462w(0) <= x_prenodeone_5_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3468w(0) <= x_prenodeone_5_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4256w(0) <= x_prenodeone_6_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4315w(0) <= x_prenodeone_6_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4321w(0) <= x_prenodeone_6_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4327w(0) <= x_prenodeone_6_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4333w(0) <= x_prenodeone_6_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4339w(0) <= x_prenodeone_6_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4345w(0) <= x_prenodeone_6_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4351w(0) <= x_prenodeone_6_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4357w(0) <= x_prenodeone_6_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4363w(0) <= x_prenodeone_6_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4369w(0) <= x_prenodeone_6_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4261w(0) <= x_prenodeone_6_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4375w(0) <= x_prenodeone_6_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4381w(0) <= x_prenodeone_6_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4387w(0) <= x_prenodeone_6_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4393w(0) <= x_prenodeone_6_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4399w(0) <= x_prenodeone_6_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4405w(0) <= x_prenodeone_6_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4411w(0) <= x_prenodeone_6_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4417w(0) <= x_prenodeone_6_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4421w(0) <= x_prenodeone_6_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4225w(0) <= x_prenodeone_6_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4267w(0) <= x_prenodeone_6_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4230w(0) <= x_prenodeone_6_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4232w(0) <= x_prenodeone_6_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4234w(0) <= x_prenodeone_6_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4236w(0) <= x_prenodeone_6_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4273w(0) <= x_prenodeone_6_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4279w(0) <= x_prenodeone_6_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4285w(0) <= x_prenodeone_6_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4291w(0) <= x_prenodeone_6_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4297w(0) <= x_prenodeone_6_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4303w(0) <= x_prenodeone_6_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4309w(0) <= x_prenodeone_6_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5092w(0) <= x_prenodeone_7_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5151w(0) <= x_prenodeone_7_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5157w(0) <= x_prenodeone_7_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5163w(0) <= x_prenodeone_7_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5169w(0) <= x_prenodeone_7_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5175w(0) <= x_prenodeone_7_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5181w(0) <= x_prenodeone_7_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5187w(0) <= x_prenodeone_7_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5193w(0) <= x_prenodeone_7_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5199w(0) <= x_prenodeone_7_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5205w(0) <= x_prenodeone_7_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5097w(0) <= x_prenodeone_7_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5211w(0) <= x_prenodeone_7_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5217w(0) <= x_prenodeone_7_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5223w(0) <= x_prenodeone_7_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5229w(0) <= x_prenodeone_7_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5235w(0) <= x_prenodeone_7_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5241w(0) <= x_prenodeone_7_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5247w(0) <= x_prenodeone_7_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5251w(0) <= x_prenodeone_7_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5057w(0) <= x_prenodeone_7_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5062w(0) <= x_prenodeone_7_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5103w(0) <= x_prenodeone_7_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5064w(0) <= x_prenodeone_7_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5066w(0) <= x_prenodeone_7_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5068w(0) <= x_prenodeone_7_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5070w(0) <= x_prenodeone_7_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5109w(0) <= x_prenodeone_7_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5115w(0) <= x_prenodeone_7_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5121w(0) <= x_prenodeone_7_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5127w(0) <= x_prenodeone_7_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5133w(0) <= x_prenodeone_7_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5139w(0) <= x_prenodeone_7_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range5145w(0) <= x_prenodeone_7_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5923w(0) <= x_prenodeone_8_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5982w(0) <= x_prenodeone_8_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5988w(0) <= x_prenodeone_8_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5994w(0) <= x_prenodeone_8_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6000w(0) <= x_prenodeone_8_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6006w(0) <= x_prenodeone_8_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6012w(0) <= x_prenodeone_8_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6018w(0) <= x_prenodeone_8_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6024w(0) <= x_prenodeone_8_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6030w(0) <= x_prenodeone_8_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6036w(0) <= x_prenodeone_8_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5928w(0) <= x_prenodeone_8_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6042w(0) <= x_prenodeone_8_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6048w(0) <= x_prenodeone_8_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6054w(0) <= x_prenodeone_8_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6060w(0) <= x_prenodeone_8_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6066w(0) <= x_prenodeone_8_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6072w(0) <= x_prenodeone_8_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range6076w(0) <= x_prenodeone_8_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5884w(0) <= x_prenodeone_8_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5889w(0) <= x_prenodeone_8_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5891w(0) <= x_prenodeone_8_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5934w(0) <= x_prenodeone_8_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5893w(0) <= x_prenodeone_8_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5895w(0) <= x_prenodeone_8_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5897w(0) <= x_prenodeone_8_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5899w(0) <= x_prenodeone_8_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5940w(0) <= x_prenodeone_8_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5946w(0) <= x_prenodeone_8_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5952w(0) <= x_prenodeone_8_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5958w(0) <= x_prenodeone_8_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5964w(0) <= x_prenodeone_8_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5970w(0) <= x_prenodeone_8_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5976w(0) <= x_prenodeone_8_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6749w(0) <= x_prenodeone_9_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6808w(0) <= x_prenodeone_9_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6814w(0) <= x_prenodeone_9_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6820w(0) <= x_prenodeone_9_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6826w(0) <= x_prenodeone_9_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6832w(0) <= x_prenodeone_9_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6838w(0) <= x_prenodeone_9_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6844w(0) <= x_prenodeone_9_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6850w(0) <= x_prenodeone_9_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6856w(0) <= x_prenodeone_9_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6862w(0) <= x_prenodeone_9_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6754w(0) <= x_prenodeone_9_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6868w(0) <= x_prenodeone_9_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6874w(0) <= x_prenodeone_9_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6880w(0) <= x_prenodeone_9_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6886w(0) <= x_prenodeone_9_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6892w(0) <= x_prenodeone_9_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6896w(0) <= x_prenodeone_9_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6706w(0) <= x_prenodeone_9_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6711w(0) <= x_prenodeone_9_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6713w(0) <= x_prenodeone_9_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6715w(0) <= x_prenodeone_9_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6760w(0) <= x_prenodeone_9_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6717w(0) <= x_prenodeone_9_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6719w(0) <= x_prenodeone_9_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6721w(0) <= x_prenodeone_9_w(32);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6723w(0) <= x_prenodeone_9_w(33);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6766w(0) <= x_prenodeone_9_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6772w(0) <= x_prenodeone_9_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6778w(0) <= x_prenodeone_9_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6784w(0) <= x_prenodeone_9_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6790w(0) <= x_prenodeone_9_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6796w(0) <= x_prenodeone_9_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6802w(0) <= x_prenodeone_9_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7714w(0) <= x_prenodetwo_10_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7743w(0) <= x_prenodetwo_10_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7746w(0) <= x_prenodetwo_10_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7749w(0) <= x_prenodetwo_10_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7752w(0) <= x_prenodetwo_10_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7755w(0) <= x_prenodetwo_10_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7758w(0) <= x_prenodetwo_10_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7761w(0) <= x_prenodetwo_10_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7764w(0) <= x_prenodetwo_10_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7767w(0) <= x_prenodetwo_10_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7770w(0) <= x_prenodetwo_10_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7716w(0) <= x_prenodetwo_10_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7773w(0) <= x_prenodetwo_10_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7776w(0) <= x_prenodetwo_10_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7779w(0) <= x_prenodetwo_10_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7544w(0) <= x_prenodetwo_10_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7548w(0) <= x_prenodetwo_10_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7550w(0) <= x_prenodetwo_10_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7552w(0) <= x_prenodetwo_10_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7554w(0) <= x_prenodetwo_10_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7556w(0) <= x_prenodetwo_10_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7558w(0) <= x_prenodetwo_10_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7719w(0) <= x_prenodetwo_10_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7560w(0) <= x_prenodetwo_10_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7562w(0) <= x_prenodetwo_10_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7564w(0) <= x_prenodetwo_10_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7566w(0) <= x_prenodetwo_10_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7722w(0) <= x_prenodetwo_10_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7725w(0) <= x_prenodetwo_10_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7728w(0) <= x_prenodetwo_10_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7731w(0) <= x_prenodetwo_10_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7734w(0) <= x_prenodetwo_10_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7737w(0) <= x_prenodetwo_10_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7740w(0) <= x_prenodetwo_10_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8524w(0) <= x_prenodetwo_11_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8553w(0) <= x_prenodetwo_11_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8556w(0) <= x_prenodetwo_11_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8559w(0) <= x_prenodetwo_11_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8562w(0) <= x_prenodetwo_11_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8565w(0) <= x_prenodetwo_11_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8568w(0) <= x_prenodetwo_11_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8571w(0) <= x_prenodetwo_11_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8574w(0) <= x_prenodetwo_11_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8577w(0) <= x_prenodetwo_11_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8580w(0) <= x_prenodetwo_11_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8526w(0) <= x_prenodetwo_11_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8583w(0) <= x_prenodetwo_11_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8586w(0) <= x_prenodetwo_11_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8358w(0) <= x_prenodetwo_11_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8362w(0) <= x_prenodetwo_11_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8364w(0) <= x_prenodetwo_11_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8366w(0) <= x_prenodetwo_11_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8368w(0) <= x_prenodetwo_11_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8370w(0) <= x_prenodetwo_11_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8372w(0) <= x_prenodetwo_11_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8374w(0) <= x_prenodetwo_11_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8529w(0) <= x_prenodetwo_11_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8376w(0) <= x_prenodetwo_11_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8378w(0) <= x_prenodetwo_11_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8380w(0) <= x_prenodetwo_11_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8382w(0) <= x_prenodetwo_11_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8532w(0) <= x_prenodetwo_11_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8535w(0) <= x_prenodetwo_11_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8538w(0) <= x_prenodetwo_11_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8541w(0) <= x_prenodetwo_11_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8544w(0) <= x_prenodetwo_11_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8547w(0) <= x_prenodetwo_11_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range8550w(0) <= x_prenodetwo_11_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9329w(0) <= x_prenodetwo_12_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9358w(0) <= x_prenodetwo_12_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9361w(0) <= x_prenodetwo_12_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9364w(0) <= x_prenodetwo_12_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9367w(0) <= x_prenodetwo_12_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9370w(0) <= x_prenodetwo_12_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9373w(0) <= x_prenodetwo_12_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9376w(0) <= x_prenodetwo_12_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9379w(0) <= x_prenodetwo_12_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9382w(0) <= x_prenodetwo_12_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9385w(0) <= x_prenodetwo_12_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9331w(0) <= x_prenodetwo_12_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9388w(0) <= x_prenodetwo_12_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9167w(0) <= x_prenodetwo_12_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9171w(0) <= x_prenodetwo_12_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9173w(0) <= x_prenodetwo_12_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9175w(0) <= x_prenodetwo_12_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9177w(0) <= x_prenodetwo_12_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9179w(0) <= x_prenodetwo_12_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9181w(0) <= x_prenodetwo_12_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9183w(0) <= x_prenodetwo_12_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9185w(0) <= x_prenodetwo_12_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9334w(0) <= x_prenodetwo_12_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9187w(0) <= x_prenodetwo_12_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9189w(0) <= x_prenodetwo_12_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9191w(0) <= x_prenodetwo_12_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9193w(0) <= x_prenodetwo_12_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9337w(0) <= x_prenodetwo_12_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9340w(0) <= x_prenodetwo_12_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9343w(0) <= x_prenodetwo_12_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9346w(0) <= x_prenodetwo_12_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9349w(0) <= x_prenodetwo_12_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9352w(0) <= x_prenodetwo_12_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range9355w(0) <= x_prenodetwo_12_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10129w(0) <= x_prenodetwo_13_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10158w(0) <= x_prenodetwo_13_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10161w(0) <= x_prenodetwo_13_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10164w(0) <= x_prenodetwo_13_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10167w(0) <= x_prenodetwo_13_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10170w(0) <= x_prenodetwo_13_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10173w(0) <= x_prenodetwo_13_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10176w(0) <= x_prenodetwo_13_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10179w(0) <= x_prenodetwo_13_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10182w(0) <= x_prenodetwo_13_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10185w(0) <= x_prenodetwo_13_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10131w(0) <= x_prenodetwo_13_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9971w(0) <= x_prenodetwo_13_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9975w(0) <= x_prenodetwo_13_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9977w(0) <= x_prenodetwo_13_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9979w(0) <= x_prenodetwo_13_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9981w(0) <= x_prenodetwo_13_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9983w(0) <= x_prenodetwo_13_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9985w(0) <= x_prenodetwo_13_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9987w(0) <= x_prenodetwo_13_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9989w(0) <= x_prenodetwo_13_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9991w(0) <= x_prenodetwo_13_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10134w(0) <= x_prenodetwo_13_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9993w(0) <= x_prenodetwo_13_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9995w(0) <= x_prenodetwo_13_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9997w(0) <= x_prenodetwo_13_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9999w(0) <= x_prenodetwo_13_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10137w(0) <= x_prenodetwo_13_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10140w(0) <= x_prenodetwo_13_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10143w(0) <= x_prenodetwo_13_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10146w(0) <= x_prenodetwo_13_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10149w(0) <= x_prenodetwo_13_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10152w(0) <= x_prenodetwo_13_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range10155w(0) <= x_prenodetwo_13_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1054w(0) <= x_prenodetwo_2_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1083w(0) <= x_prenodetwo_2_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1086w(0) <= x_prenodetwo_2_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1089w(0) <= x_prenodetwo_2_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1092w(0) <= x_prenodetwo_2_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1095w(0) <= x_prenodetwo_2_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1098w(0) <= x_prenodetwo_2_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1101w(0) <= x_prenodetwo_2_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1104w(0) <= x_prenodetwo_2_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1107w(0) <= x_prenodetwo_2_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1110w(0) <= x_prenodetwo_2_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1056w(0) <= x_prenodetwo_2_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1113w(0) <= x_prenodetwo_2_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1116w(0) <= x_prenodetwo_2_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1119w(0) <= x_prenodetwo_2_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1122w(0) <= x_prenodetwo_2_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1125w(0) <= x_prenodetwo_2_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1128w(0) <= x_prenodetwo_2_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1131w(0) <= x_prenodetwo_2_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1134w(0) <= x_prenodetwo_2_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1137w(0) <= x_prenodetwo_2_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1140w(0) <= x_prenodetwo_2_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1059w(0) <= x_prenodetwo_2_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1143w(0) <= x_prenodetwo_2_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range852w(0) <= x_prenodetwo_2_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range856w(0) <= x_prenodetwo_2_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range858w(0) <= x_prenodetwo_2_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1062w(0) <= x_prenodetwo_2_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1065w(0) <= x_prenodetwo_2_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1068w(0) <= x_prenodetwo_2_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1071w(0) <= x_prenodetwo_2_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1074w(0) <= x_prenodetwo_2_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1077w(0) <= x_prenodetwo_2_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range1080w(0) <= x_prenodetwo_2_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1904w(0) <= x_prenodetwo_3_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1933w(0) <= x_prenodetwo_3_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1936w(0) <= x_prenodetwo_3_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1939w(0) <= x_prenodetwo_3_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1942w(0) <= x_prenodetwo_3_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1945w(0) <= x_prenodetwo_3_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1948w(0) <= x_prenodetwo_3_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1951w(0) <= x_prenodetwo_3_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1954w(0) <= x_prenodetwo_3_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1957w(0) <= x_prenodetwo_3_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1960w(0) <= x_prenodetwo_3_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1906w(0) <= x_prenodetwo_3_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1963w(0) <= x_prenodetwo_3_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1966w(0) <= x_prenodetwo_3_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1969w(0) <= x_prenodetwo_3_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1972w(0) <= x_prenodetwo_3_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1975w(0) <= x_prenodetwo_3_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1978w(0) <= x_prenodetwo_3_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1981w(0) <= x_prenodetwo_3_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1984w(0) <= x_prenodetwo_3_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1987w(0) <= x_prenodetwo_3_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1990w(0) <= x_prenodetwo_3_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1909w(0) <= x_prenodetwo_3_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1706w(0) <= x_prenodetwo_3_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1710w(0) <= x_prenodetwo_3_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1712w(0) <= x_prenodetwo_3_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1714w(0) <= x_prenodetwo_3_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1912w(0) <= x_prenodetwo_3_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1915w(0) <= x_prenodetwo_3_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1918w(0) <= x_prenodetwo_3_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1921w(0) <= x_prenodetwo_3_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1924w(0) <= x_prenodetwo_3_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1927w(0) <= x_prenodetwo_3_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1930w(0) <= x_prenodetwo_3_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2749w(0) <= x_prenodetwo_4_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2778w(0) <= x_prenodetwo_4_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2781w(0) <= x_prenodetwo_4_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2784w(0) <= x_prenodetwo_4_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2787w(0) <= x_prenodetwo_4_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2790w(0) <= x_prenodetwo_4_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2793w(0) <= x_prenodetwo_4_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2796w(0) <= x_prenodetwo_4_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2799w(0) <= x_prenodetwo_4_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2802w(0) <= x_prenodetwo_4_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2805w(0) <= x_prenodetwo_4_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2751w(0) <= x_prenodetwo_4_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2808w(0) <= x_prenodetwo_4_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2811w(0) <= x_prenodetwo_4_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2814w(0) <= x_prenodetwo_4_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2817w(0) <= x_prenodetwo_4_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2820w(0) <= x_prenodetwo_4_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2823w(0) <= x_prenodetwo_4_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2826w(0) <= x_prenodetwo_4_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2829w(0) <= x_prenodetwo_4_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2832w(0) <= x_prenodetwo_4_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2555w(0) <= x_prenodetwo_4_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2754w(0) <= x_prenodetwo_4_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2559w(0) <= x_prenodetwo_4_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2561w(0) <= x_prenodetwo_4_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2563w(0) <= x_prenodetwo_4_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2565w(0) <= x_prenodetwo_4_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2757w(0) <= x_prenodetwo_4_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2760w(0) <= x_prenodetwo_4_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2763w(0) <= x_prenodetwo_4_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2766w(0) <= x_prenodetwo_4_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2769w(0) <= x_prenodetwo_4_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2772w(0) <= x_prenodetwo_4_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2775w(0) <= x_prenodetwo_4_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3589w(0) <= x_prenodetwo_5_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3618w(0) <= x_prenodetwo_5_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3621w(0) <= x_prenodetwo_5_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3624w(0) <= x_prenodetwo_5_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3627w(0) <= x_prenodetwo_5_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3630w(0) <= x_prenodetwo_5_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3633w(0) <= x_prenodetwo_5_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3636w(0) <= x_prenodetwo_5_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3639w(0) <= x_prenodetwo_5_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3642w(0) <= x_prenodetwo_5_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3645w(0) <= x_prenodetwo_5_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3591w(0) <= x_prenodetwo_5_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3648w(0) <= x_prenodetwo_5_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3651w(0) <= x_prenodetwo_5_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3654w(0) <= x_prenodetwo_5_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3657w(0) <= x_prenodetwo_5_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3660w(0) <= x_prenodetwo_5_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3663w(0) <= x_prenodetwo_5_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3666w(0) <= x_prenodetwo_5_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3669w(0) <= x_prenodetwo_5_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3399w(0) <= x_prenodetwo_5_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3403w(0) <= x_prenodetwo_5_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3594w(0) <= x_prenodetwo_5_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3405w(0) <= x_prenodetwo_5_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3407w(0) <= x_prenodetwo_5_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3409w(0) <= x_prenodetwo_5_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3411w(0) <= x_prenodetwo_5_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3597w(0) <= x_prenodetwo_5_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3600w(0) <= x_prenodetwo_5_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3603w(0) <= x_prenodetwo_5_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3606w(0) <= x_prenodetwo_5_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3609w(0) <= x_prenodetwo_5_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3612w(0) <= x_prenodetwo_5_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3615w(0) <= x_prenodetwo_5_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4424w(0) <= x_prenodetwo_6_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4453w(0) <= x_prenodetwo_6_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4456w(0) <= x_prenodetwo_6_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4459w(0) <= x_prenodetwo_6_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4462w(0) <= x_prenodetwo_6_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4465w(0) <= x_prenodetwo_6_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4468w(0) <= x_prenodetwo_6_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4471w(0) <= x_prenodetwo_6_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4474w(0) <= x_prenodetwo_6_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4477w(0) <= x_prenodetwo_6_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4480w(0) <= x_prenodetwo_6_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4426w(0) <= x_prenodetwo_6_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4483w(0) <= x_prenodetwo_6_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4486w(0) <= x_prenodetwo_6_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4489w(0) <= x_prenodetwo_6_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4492w(0) <= x_prenodetwo_6_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4495w(0) <= x_prenodetwo_6_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4498w(0) <= x_prenodetwo_6_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4501w(0) <= x_prenodetwo_6_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4238w(0) <= x_prenodetwo_6_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4242w(0) <= x_prenodetwo_6_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4244w(0) <= x_prenodetwo_6_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4429w(0) <= x_prenodetwo_6_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4246w(0) <= x_prenodetwo_6_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4248w(0) <= x_prenodetwo_6_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4250w(0) <= x_prenodetwo_6_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4252w(0) <= x_prenodetwo_6_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4432w(0) <= x_prenodetwo_6_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4435w(0) <= x_prenodetwo_6_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4438w(0) <= x_prenodetwo_6_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4441w(0) <= x_prenodetwo_6_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4444w(0) <= x_prenodetwo_6_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4447w(0) <= x_prenodetwo_6_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4450w(0) <= x_prenodetwo_6_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5254w(0) <= x_prenodetwo_7_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5283w(0) <= x_prenodetwo_7_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5286w(0) <= x_prenodetwo_7_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5289w(0) <= x_prenodetwo_7_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5292w(0) <= x_prenodetwo_7_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5295w(0) <= x_prenodetwo_7_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5298w(0) <= x_prenodetwo_7_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5301w(0) <= x_prenodetwo_7_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5304w(0) <= x_prenodetwo_7_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5307w(0) <= x_prenodetwo_7_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5310w(0) <= x_prenodetwo_7_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5256w(0) <= x_prenodetwo_7_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5313w(0) <= x_prenodetwo_7_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5316w(0) <= x_prenodetwo_7_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5319w(0) <= x_prenodetwo_7_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5322w(0) <= x_prenodetwo_7_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5325w(0) <= x_prenodetwo_7_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5328w(0) <= x_prenodetwo_7_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5072w(0) <= x_prenodetwo_7_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5076w(0) <= x_prenodetwo_7_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5078w(0) <= x_prenodetwo_7_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5080w(0) <= x_prenodetwo_7_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5259w(0) <= x_prenodetwo_7_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5082w(0) <= x_prenodetwo_7_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5084w(0) <= x_prenodetwo_7_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5086w(0) <= x_prenodetwo_7_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5088w(0) <= x_prenodetwo_7_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5262w(0) <= x_prenodetwo_7_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5265w(0) <= x_prenodetwo_7_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5268w(0) <= x_prenodetwo_7_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5271w(0) <= x_prenodetwo_7_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5274w(0) <= x_prenodetwo_7_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5277w(0) <= x_prenodetwo_7_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range5280w(0) <= x_prenodetwo_7_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6079w(0) <= x_prenodetwo_8_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6108w(0) <= x_prenodetwo_8_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6111w(0) <= x_prenodetwo_8_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6114w(0) <= x_prenodetwo_8_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6117w(0) <= x_prenodetwo_8_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6120w(0) <= x_prenodetwo_8_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6123w(0) <= x_prenodetwo_8_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6126w(0) <= x_prenodetwo_8_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6129w(0) <= x_prenodetwo_8_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6132w(0) <= x_prenodetwo_8_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6135w(0) <= x_prenodetwo_8_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6081w(0) <= x_prenodetwo_8_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6138w(0) <= x_prenodetwo_8_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6141w(0) <= x_prenodetwo_8_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6144w(0) <= x_prenodetwo_8_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6147w(0) <= x_prenodetwo_8_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6150w(0) <= x_prenodetwo_8_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5901w(0) <= x_prenodetwo_8_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5905w(0) <= x_prenodetwo_8_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5907w(0) <= x_prenodetwo_8_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5909w(0) <= x_prenodetwo_8_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5911w(0) <= x_prenodetwo_8_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6084w(0) <= x_prenodetwo_8_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5913w(0) <= x_prenodetwo_8_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5915w(0) <= x_prenodetwo_8_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5917w(0) <= x_prenodetwo_8_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5919w(0) <= x_prenodetwo_8_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6087w(0) <= x_prenodetwo_8_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6090w(0) <= x_prenodetwo_8_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6093w(0) <= x_prenodetwo_8_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6096w(0) <= x_prenodetwo_8_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6099w(0) <= x_prenodetwo_8_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6102w(0) <= x_prenodetwo_8_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range6105w(0) <= x_prenodetwo_8_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6899w(0) <= x_prenodetwo_9_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6928w(0) <= x_prenodetwo_9_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6931w(0) <= x_prenodetwo_9_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6934w(0) <= x_prenodetwo_9_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6937w(0) <= x_prenodetwo_9_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6940w(0) <= x_prenodetwo_9_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6943w(0) <= x_prenodetwo_9_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6946w(0) <= x_prenodetwo_9_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6949w(0) <= x_prenodetwo_9_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6952w(0) <= x_prenodetwo_9_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6955w(0) <= x_prenodetwo_9_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6901w(0) <= x_prenodetwo_9_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6958w(0) <= x_prenodetwo_9_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6961w(0) <= x_prenodetwo_9_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6964w(0) <= x_prenodetwo_9_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6967w(0) <= x_prenodetwo_9_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6725w(0) <= x_prenodetwo_9_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6729w(0) <= x_prenodetwo_9_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6731w(0) <= x_prenodetwo_9_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6733w(0) <= x_prenodetwo_9_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6735w(0) <= x_prenodetwo_9_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6737w(0) <= x_prenodetwo_9_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6904w(0) <= x_prenodetwo_9_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6739w(0) <= x_prenodetwo_9_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6741w(0) <= x_prenodetwo_9_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6743w(0) <= x_prenodetwo_9_w(32);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6745w(0) <= x_prenodetwo_9_w(33);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6907w(0) <= x_prenodetwo_9_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6910w(0) <= x_prenodetwo_9_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6913w(0) <= x_prenodetwo_9_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6916w(0) <= x_prenodetwo_9_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6919w(0) <= x_prenodetwo_9_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6922w(0) <= x_prenodetwo_9_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6925w(0) <= x_prenodetwo_9_w(9);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7791w(0) <= y_prenode_10_w(0);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7872w(0) <= y_prenode_10_w(10);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7880w(0) <= y_prenode_10_w(11);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7888w(0) <= y_prenode_10_w(12);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7896w(0) <= y_prenode_10_w(13);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7904w(0) <= y_prenode_10_w(14);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7912w(0) <= y_prenode_10_w(15);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7920w(0) <= y_prenode_10_w(16);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7928w(0) <= y_prenode_10_w(17);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7936w(0) <= y_prenode_10_w(18);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7944w(0) <= y_prenode_10_w(19);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7800w(0) <= y_prenode_10_w(1);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7952w(0) <= y_prenode_10_w(20);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7960w(0) <= y_prenode_10_w(21);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7968w(0) <= y_prenode_10_w(22);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7976w(0) <= y_prenode_10_w(23);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7984w(0) <= y_prenode_10_w(24);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7992w(0) <= y_prenode_10_w(25);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8000w(0) <= y_prenode_10_w(26);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8008w(0) <= y_prenode_10_w(27);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8016w(0) <= y_prenode_10_w(28);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8024w(0) <= y_prenode_10_w(29);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7808w(0) <= y_prenode_10_w(2);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8032w(0) <= y_prenode_10_w(30);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8040w(0) <= y_prenode_10_w(31);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8048w(0) <= y_prenode_10_w(32);
	wire_ccc_cordic_m_w_y_prenode_10_w_range8056w(0) <= y_prenode_10_w(33);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7816w(0) <= y_prenode_10_w(3);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7824w(0) <= y_prenode_10_w(4);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7832w(0) <= y_prenode_10_w(5);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7840w(0) <= y_prenode_10_w(6);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7848w(0) <= y_prenode_10_w(7);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7856w(0) <= y_prenode_10_w(8);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7864w(0) <= y_prenode_10_w(9);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8598w(0) <= y_prenode_11_w(0);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8679w(0) <= y_prenode_11_w(10);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8687w(0) <= y_prenode_11_w(11);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8695w(0) <= y_prenode_11_w(12);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8703w(0) <= y_prenode_11_w(13);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8711w(0) <= y_prenode_11_w(14);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8719w(0) <= y_prenode_11_w(15);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8727w(0) <= y_prenode_11_w(16);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8735w(0) <= y_prenode_11_w(17);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8743w(0) <= y_prenode_11_w(18);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8751w(0) <= y_prenode_11_w(19);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8607w(0) <= y_prenode_11_w(1);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8759w(0) <= y_prenode_11_w(20);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8767w(0) <= y_prenode_11_w(21);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8775w(0) <= y_prenode_11_w(22);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8783w(0) <= y_prenode_11_w(23);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8791w(0) <= y_prenode_11_w(24);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8799w(0) <= y_prenode_11_w(25);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8807w(0) <= y_prenode_11_w(26);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8815w(0) <= y_prenode_11_w(27);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8823w(0) <= y_prenode_11_w(28);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8831w(0) <= y_prenode_11_w(29);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8615w(0) <= y_prenode_11_w(2);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8839w(0) <= y_prenode_11_w(30);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8847w(0) <= y_prenode_11_w(31);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8855w(0) <= y_prenode_11_w(32);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8863w(0) <= y_prenode_11_w(33);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8623w(0) <= y_prenode_11_w(3);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8631w(0) <= y_prenode_11_w(4);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8639w(0) <= y_prenode_11_w(5);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8647w(0) <= y_prenode_11_w(6);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8655w(0) <= y_prenode_11_w(7);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8663w(0) <= y_prenode_11_w(8);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8671w(0) <= y_prenode_11_w(9);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9400w(0) <= y_prenode_12_w(0);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9481w(0) <= y_prenode_12_w(10);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9489w(0) <= y_prenode_12_w(11);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9497w(0) <= y_prenode_12_w(12);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9505w(0) <= y_prenode_12_w(13);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9513w(0) <= y_prenode_12_w(14);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9521w(0) <= y_prenode_12_w(15);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9529w(0) <= y_prenode_12_w(16);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9537w(0) <= y_prenode_12_w(17);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9545w(0) <= y_prenode_12_w(18);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9553w(0) <= y_prenode_12_w(19);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9409w(0) <= y_prenode_12_w(1);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9561w(0) <= y_prenode_12_w(20);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9569w(0) <= y_prenode_12_w(21);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9577w(0) <= y_prenode_12_w(22);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9585w(0) <= y_prenode_12_w(23);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9593w(0) <= y_prenode_12_w(24);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9601w(0) <= y_prenode_12_w(25);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9609w(0) <= y_prenode_12_w(26);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9617w(0) <= y_prenode_12_w(27);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9625w(0) <= y_prenode_12_w(28);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9633w(0) <= y_prenode_12_w(29);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9417w(0) <= y_prenode_12_w(2);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9641w(0) <= y_prenode_12_w(30);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9649w(0) <= y_prenode_12_w(31);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9657w(0) <= y_prenode_12_w(32);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9665w(0) <= y_prenode_12_w(33);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9425w(0) <= y_prenode_12_w(3);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9433w(0) <= y_prenode_12_w(4);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9441w(0) <= y_prenode_12_w(5);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9449w(0) <= y_prenode_12_w(6);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9457w(0) <= y_prenode_12_w(7);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9465w(0) <= y_prenode_12_w(8);
	wire_ccc_cordic_m_w_y_prenode_12_w_range9473w(0) <= y_prenode_12_w(9);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10197w(0) <= y_prenode_13_w(0);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10278w(0) <= y_prenode_13_w(10);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10286w(0) <= y_prenode_13_w(11);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10294w(0) <= y_prenode_13_w(12);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10302w(0) <= y_prenode_13_w(13);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10310w(0) <= y_prenode_13_w(14);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10318w(0) <= y_prenode_13_w(15);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10326w(0) <= y_prenode_13_w(16);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10334w(0) <= y_prenode_13_w(17);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10342w(0) <= y_prenode_13_w(18);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10350w(0) <= y_prenode_13_w(19);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10206w(0) <= y_prenode_13_w(1);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10358w(0) <= y_prenode_13_w(20);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10366w(0) <= y_prenode_13_w(21);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10374w(0) <= y_prenode_13_w(22);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10382w(0) <= y_prenode_13_w(23);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10390w(0) <= y_prenode_13_w(24);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10398w(0) <= y_prenode_13_w(25);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10406w(0) <= y_prenode_13_w(26);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10414w(0) <= y_prenode_13_w(27);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10422w(0) <= y_prenode_13_w(28);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10430w(0) <= y_prenode_13_w(29);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10214w(0) <= y_prenode_13_w(2);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10438w(0) <= y_prenode_13_w(30);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10446w(0) <= y_prenode_13_w(31);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10454w(0) <= y_prenode_13_w(32);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10462w(0) <= y_prenode_13_w(33);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10222w(0) <= y_prenode_13_w(3);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10230w(0) <= y_prenode_13_w(4);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10238w(0) <= y_prenode_13_w(5);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10246w(0) <= y_prenode_13_w(6);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10254w(0) <= y_prenode_13_w(7);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10262w(0) <= y_prenode_13_w(8);
	wire_ccc_cordic_m_w_y_prenode_13_w_range10270w(0) <= y_prenode_13_w(9);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1155w(0) <= y_prenode_2_w(0);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1236w(0) <= y_prenode_2_w(10);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1244w(0) <= y_prenode_2_w(11);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1252w(0) <= y_prenode_2_w(12);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1260w(0) <= y_prenode_2_w(13);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1268w(0) <= y_prenode_2_w(14);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1276w(0) <= y_prenode_2_w(15);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1284w(0) <= y_prenode_2_w(16);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1292w(0) <= y_prenode_2_w(17);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1300w(0) <= y_prenode_2_w(18);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1308w(0) <= y_prenode_2_w(19);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1164w(0) <= y_prenode_2_w(1);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1316w(0) <= y_prenode_2_w(20);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1324w(0) <= y_prenode_2_w(21);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1332w(0) <= y_prenode_2_w(22);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1340w(0) <= y_prenode_2_w(23);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1348w(0) <= y_prenode_2_w(24);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1356w(0) <= y_prenode_2_w(25);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1364w(0) <= y_prenode_2_w(26);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1372w(0) <= y_prenode_2_w(27);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1380w(0) <= y_prenode_2_w(28);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1388w(0) <= y_prenode_2_w(29);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1172w(0) <= y_prenode_2_w(2);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1396w(0) <= y_prenode_2_w(30);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1404w(0) <= y_prenode_2_w(31);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1412w(0) <= y_prenode_2_w(32);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1420w(0) <= y_prenode_2_w(33);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1180w(0) <= y_prenode_2_w(3);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1188w(0) <= y_prenode_2_w(4);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1196w(0) <= y_prenode_2_w(5);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1204w(0) <= y_prenode_2_w(6);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1212w(0) <= y_prenode_2_w(7);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1220w(0) <= y_prenode_2_w(8);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1228w(0) <= y_prenode_2_w(9);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2002w(0) <= y_prenode_3_w(0);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2083w(0) <= y_prenode_3_w(10);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2091w(0) <= y_prenode_3_w(11);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2099w(0) <= y_prenode_3_w(12);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2107w(0) <= y_prenode_3_w(13);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2115w(0) <= y_prenode_3_w(14);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2123w(0) <= y_prenode_3_w(15);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2131w(0) <= y_prenode_3_w(16);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2139w(0) <= y_prenode_3_w(17);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2147w(0) <= y_prenode_3_w(18);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2155w(0) <= y_prenode_3_w(19);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2011w(0) <= y_prenode_3_w(1);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2163w(0) <= y_prenode_3_w(20);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2171w(0) <= y_prenode_3_w(21);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2179w(0) <= y_prenode_3_w(22);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2187w(0) <= y_prenode_3_w(23);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2195w(0) <= y_prenode_3_w(24);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2203w(0) <= y_prenode_3_w(25);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2211w(0) <= y_prenode_3_w(26);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2219w(0) <= y_prenode_3_w(27);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2227w(0) <= y_prenode_3_w(28);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2235w(0) <= y_prenode_3_w(29);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2019w(0) <= y_prenode_3_w(2);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2243w(0) <= y_prenode_3_w(30);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2251w(0) <= y_prenode_3_w(31);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2259w(0) <= y_prenode_3_w(32);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2267w(0) <= y_prenode_3_w(33);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2027w(0) <= y_prenode_3_w(3);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2035w(0) <= y_prenode_3_w(4);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2043w(0) <= y_prenode_3_w(5);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2051w(0) <= y_prenode_3_w(6);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2059w(0) <= y_prenode_3_w(7);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2067w(0) <= y_prenode_3_w(8);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2075w(0) <= y_prenode_3_w(9);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2844w(0) <= y_prenode_4_w(0);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2925w(0) <= y_prenode_4_w(10);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2933w(0) <= y_prenode_4_w(11);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2941w(0) <= y_prenode_4_w(12);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2949w(0) <= y_prenode_4_w(13);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2957w(0) <= y_prenode_4_w(14);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2965w(0) <= y_prenode_4_w(15);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2973w(0) <= y_prenode_4_w(16);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2981w(0) <= y_prenode_4_w(17);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2989w(0) <= y_prenode_4_w(18);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2997w(0) <= y_prenode_4_w(19);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2853w(0) <= y_prenode_4_w(1);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3005w(0) <= y_prenode_4_w(20);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3013w(0) <= y_prenode_4_w(21);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3021w(0) <= y_prenode_4_w(22);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3029w(0) <= y_prenode_4_w(23);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3037w(0) <= y_prenode_4_w(24);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3045w(0) <= y_prenode_4_w(25);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3053w(0) <= y_prenode_4_w(26);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3061w(0) <= y_prenode_4_w(27);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3069w(0) <= y_prenode_4_w(28);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3077w(0) <= y_prenode_4_w(29);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2861w(0) <= y_prenode_4_w(2);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3085w(0) <= y_prenode_4_w(30);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3093w(0) <= y_prenode_4_w(31);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3101w(0) <= y_prenode_4_w(32);
	wire_ccc_cordic_m_w_y_prenode_4_w_range3109w(0) <= y_prenode_4_w(33);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2869w(0) <= y_prenode_4_w(3);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2877w(0) <= y_prenode_4_w(4);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2885w(0) <= y_prenode_4_w(5);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2893w(0) <= y_prenode_4_w(6);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2901w(0) <= y_prenode_4_w(7);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2909w(0) <= y_prenode_4_w(8);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2917w(0) <= y_prenode_4_w(9);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3681w(0) <= y_prenode_5_w(0);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3762w(0) <= y_prenode_5_w(10);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3770w(0) <= y_prenode_5_w(11);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3778w(0) <= y_prenode_5_w(12);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3786w(0) <= y_prenode_5_w(13);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3794w(0) <= y_prenode_5_w(14);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3802w(0) <= y_prenode_5_w(15);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3810w(0) <= y_prenode_5_w(16);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3818w(0) <= y_prenode_5_w(17);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3826w(0) <= y_prenode_5_w(18);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3834w(0) <= y_prenode_5_w(19);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3690w(0) <= y_prenode_5_w(1);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3842w(0) <= y_prenode_5_w(20);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3850w(0) <= y_prenode_5_w(21);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3858w(0) <= y_prenode_5_w(22);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3866w(0) <= y_prenode_5_w(23);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3874w(0) <= y_prenode_5_w(24);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3882w(0) <= y_prenode_5_w(25);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3890w(0) <= y_prenode_5_w(26);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3898w(0) <= y_prenode_5_w(27);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3906w(0) <= y_prenode_5_w(28);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3914w(0) <= y_prenode_5_w(29);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3698w(0) <= y_prenode_5_w(2);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3922w(0) <= y_prenode_5_w(30);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3930w(0) <= y_prenode_5_w(31);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3938w(0) <= y_prenode_5_w(32);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3946w(0) <= y_prenode_5_w(33);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3706w(0) <= y_prenode_5_w(3);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3714w(0) <= y_prenode_5_w(4);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3722w(0) <= y_prenode_5_w(5);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3730w(0) <= y_prenode_5_w(6);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3738w(0) <= y_prenode_5_w(7);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3746w(0) <= y_prenode_5_w(8);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3754w(0) <= y_prenode_5_w(9);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4513w(0) <= y_prenode_6_w(0);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4594w(0) <= y_prenode_6_w(10);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4602w(0) <= y_prenode_6_w(11);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4610w(0) <= y_prenode_6_w(12);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4618w(0) <= y_prenode_6_w(13);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4626w(0) <= y_prenode_6_w(14);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4634w(0) <= y_prenode_6_w(15);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4642w(0) <= y_prenode_6_w(16);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4650w(0) <= y_prenode_6_w(17);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4658w(0) <= y_prenode_6_w(18);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4666w(0) <= y_prenode_6_w(19);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4522w(0) <= y_prenode_6_w(1);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4674w(0) <= y_prenode_6_w(20);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4682w(0) <= y_prenode_6_w(21);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4690w(0) <= y_prenode_6_w(22);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4698w(0) <= y_prenode_6_w(23);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4706w(0) <= y_prenode_6_w(24);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4714w(0) <= y_prenode_6_w(25);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4722w(0) <= y_prenode_6_w(26);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4730w(0) <= y_prenode_6_w(27);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4738w(0) <= y_prenode_6_w(28);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4746w(0) <= y_prenode_6_w(29);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4530w(0) <= y_prenode_6_w(2);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4754w(0) <= y_prenode_6_w(30);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4762w(0) <= y_prenode_6_w(31);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4770w(0) <= y_prenode_6_w(32);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4778w(0) <= y_prenode_6_w(33);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4538w(0) <= y_prenode_6_w(3);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4546w(0) <= y_prenode_6_w(4);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4554w(0) <= y_prenode_6_w(5);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4562w(0) <= y_prenode_6_w(6);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4570w(0) <= y_prenode_6_w(7);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4578w(0) <= y_prenode_6_w(8);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4586w(0) <= y_prenode_6_w(9);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5340w(0) <= y_prenode_7_w(0);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5421w(0) <= y_prenode_7_w(10);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5429w(0) <= y_prenode_7_w(11);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5437w(0) <= y_prenode_7_w(12);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5445w(0) <= y_prenode_7_w(13);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5453w(0) <= y_prenode_7_w(14);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5461w(0) <= y_prenode_7_w(15);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5469w(0) <= y_prenode_7_w(16);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5477w(0) <= y_prenode_7_w(17);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5485w(0) <= y_prenode_7_w(18);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5493w(0) <= y_prenode_7_w(19);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5349w(0) <= y_prenode_7_w(1);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5501w(0) <= y_prenode_7_w(20);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5509w(0) <= y_prenode_7_w(21);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5517w(0) <= y_prenode_7_w(22);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5525w(0) <= y_prenode_7_w(23);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5533w(0) <= y_prenode_7_w(24);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5541w(0) <= y_prenode_7_w(25);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5549w(0) <= y_prenode_7_w(26);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5557w(0) <= y_prenode_7_w(27);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5565w(0) <= y_prenode_7_w(28);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5573w(0) <= y_prenode_7_w(29);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5357w(0) <= y_prenode_7_w(2);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5581w(0) <= y_prenode_7_w(30);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5589w(0) <= y_prenode_7_w(31);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5597w(0) <= y_prenode_7_w(32);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5605w(0) <= y_prenode_7_w(33);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5365w(0) <= y_prenode_7_w(3);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5373w(0) <= y_prenode_7_w(4);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5381w(0) <= y_prenode_7_w(5);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5389w(0) <= y_prenode_7_w(6);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5397w(0) <= y_prenode_7_w(7);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5405w(0) <= y_prenode_7_w(8);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5413w(0) <= y_prenode_7_w(9);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6162w(0) <= y_prenode_8_w(0);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6243w(0) <= y_prenode_8_w(10);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6251w(0) <= y_prenode_8_w(11);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6259w(0) <= y_prenode_8_w(12);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6267w(0) <= y_prenode_8_w(13);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6275w(0) <= y_prenode_8_w(14);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6283w(0) <= y_prenode_8_w(15);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6291w(0) <= y_prenode_8_w(16);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6299w(0) <= y_prenode_8_w(17);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6307w(0) <= y_prenode_8_w(18);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6315w(0) <= y_prenode_8_w(19);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6171w(0) <= y_prenode_8_w(1);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6323w(0) <= y_prenode_8_w(20);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6331w(0) <= y_prenode_8_w(21);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6339w(0) <= y_prenode_8_w(22);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6347w(0) <= y_prenode_8_w(23);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6355w(0) <= y_prenode_8_w(24);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6363w(0) <= y_prenode_8_w(25);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6371w(0) <= y_prenode_8_w(26);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6379w(0) <= y_prenode_8_w(27);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6387w(0) <= y_prenode_8_w(28);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6395w(0) <= y_prenode_8_w(29);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6179w(0) <= y_prenode_8_w(2);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6403w(0) <= y_prenode_8_w(30);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6411w(0) <= y_prenode_8_w(31);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6419w(0) <= y_prenode_8_w(32);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6427w(0) <= y_prenode_8_w(33);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6187w(0) <= y_prenode_8_w(3);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6195w(0) <= y_prenode_8_w(4);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6203w(0) <= y_prenode_8_w(5);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6211w(0) <= y_prenode_8_w(6);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6219w(0) <= y_prenode_8_w(7);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6227w(0) <= y_prenode_8_w(8);
	wire_ccc_cordic_m_w_y_prenode_8_w_range6235w(0) <= y_prenode_8_w(9);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6979w(0) <= y_prenode_9_w(0);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7060w(0) <= y_prenode_9_w(10);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7068w(0) <= y_prenode_9_w(11);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7076w(0) <= y_prenode_9_w(12);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7084w(0) <= y_prenode_9_w(13);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7092w(0) <= y_prenode_9_w(14);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7100w(0) <= y_prenode_9_w(15);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7108w(0) <= y_prenode_9_w(16);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7116w(0) <= y_prenode_9_w(17);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7124w(0) <= y_prenode_9_w(18);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7132w(0) <= y_prenode_9_w(19);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6988w(0) <= y_prenode_9_w(1);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7140w(0) <= y_prenode_9_w(20);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7148w(0) <= y_prenode_9_w(21);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7156w(0) <= y_prenode_9_w(22);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7164w(0) <= y_prenode_9_w(23);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7172w(0) <= y_prenode_9_w(24);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7180w(0) <= y_prenode_9_w(25);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7188w(0) <= y_prenode_9_w(26);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7196w(0) <= y_prenode_9_w(27);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7204w(0) <= y_prenode_9_w(28);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7212w(0) <= y_prenode_9_w(29);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6996w(0) <= y_prenode_9_w(2);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7220w(0) <= y_prenode_9_w(30);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7228w(0) <= y_prenode_9_w(31);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7236w(0) <= y_prenode_9_w(32);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7244w(0) <= y_prenode_9_w(33);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7004w(0) <= y_prenode_9_w(3);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7012w(0) <= y_prenode_9_w(4);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7020w(0) <= y_prenode_9_w(5);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7028w(0) <= y_prenode_9_w(6);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7036w(0) <= y_prenode_9_w(7);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7044w(0) <= y_prenode_9_w(8);
	wire_ccc_cordic_m_w_y_prenode_9_w_range7052w(0) <= y_prenode_9_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7572w(0) <= y_prenodeone_10_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7631w(0) <= y_prenodeone_10_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7637w(0) <= y_prenodeone_10_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7643w(0) <= y_prenodeone_10_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7649w(0) <= y_prenodeone_10_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7655w(0) <= y_prenodeone_10_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7661w(0) <= y_prenodeone_10_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7667w(0) <= y_prenodeone_10_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7673w(0) <= y_prenodeone_10_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7679w(0) <= y_prenodeone_10_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7685w(0) <= y_prenodeone_10_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7577w(0) <= y_prenodeone_10_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7691w(0) <= y_prenodeone_10_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7697w(0) <= y_prenodeone_10_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7703w(0) <= y_prenodeone_10_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7709w(0) <= y_prenodeone_10_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7712w(0) <= y_prenodeone_10_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7526w(0) <= y_prenodeone_10_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7529w(0) <= y_prenodeone_10_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7531w(0) <= y_prenodeone_10_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7533w(0) <= y_prenodeone_10_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7535w(0) <= y_prenodeone_10_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7583w(0) <= y_prenodeone_10_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7537w(0) <= y_prenodeone_10_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7539w(0) <= y_prenodeone_10_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7541w(0) <= y_prenodeone_10_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7543w(0) <= y_prenodeone_10_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7589w(0) <= y_prenodeone_10_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7595w(0) <= y_prenodeone_10_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7601w(0) <= y_prenodeone_10_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7607w(0) <= y_prenodeone_10_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7613w(0) <= y_prenodeone_10_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7619w(0) <= y_prenodeone_10_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7625w(0) <= y_prenodeone_10_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8388w(0) <= y_prenodeone_11_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8447w(0) <= y_prenodeone_11_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8453w(0) <= y_prenodeone_11_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8459w(0) <= y_prenodeone_11_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8465w(0) <= y_prenodeone_11_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8471w(0) <= y_prenodeone_11_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8477w(0) <= y_prenodeone_11_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8483w(0) <= y_prenodeone_11_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8489w(0) <= y_prenodeone_11_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8495w(0) <= y_prenodeone_11_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8501w(0) <= y_prenodeone_11_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8393w(0) <= y_prenodeone_11_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8507w(0) <= y_prenodeone_11_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8513w(0) <= y_prenodeone_11_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8519w(0) <= y_prenodeone_11_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8522w(0) <= y_prenodeone_11_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8338w(0) <= y_prenodeone_11_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8341w(0) <= y_prenodeone_11_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8343w(0) <= y_prenodeone_11_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8345w(0) <= y_prenodeone_11_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8347w(0) <= y_prenodeone_11_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8349w(0) <= y_prenodeone_11_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8399w(0) <= y_prenodeone_11_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8351w(0) <= y_prenodeone_11_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8353w(0) <= y_prenodeone_11_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8355w(0) <= y_prenodeone_11_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8357w(0) <= y_prenodeone_11_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8405w(0) <= y_prenodeone_11_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8411w(0) <= y_prenodeone_11_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8417w(0) <= y_prenodeone_11_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8423w(0) <= y_prenodeone_11_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8429w(0) <= y_prenodeone_11_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8435w(0) <= y_prenodeone_11_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range8441w(0) <= y_prenodeone_11_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9199w(0) <= y_prenodeone_12_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9258w(0) <= y_prenodeone_12_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9264w(0) <= y_prenodeone_12_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9270w(0) <= y_prenodeone_12_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9276w(0) <= y_prenodeone_12_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9282w(0) <= y_prenodeone_12_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9288w(0) <= y_prenodeone_12_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9294w(0) <= y_prenodeone_12_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9300w(0) <= y_prenodeone_12_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9306w(0) <= y_prenodeone_12_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9312w(0) <= y_prenodeone_12_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9204w(0) <= y_prenodeone_12_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9318w(0) <= y_prenodeone_12_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9324w(0) <= y_prenodeone_12_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9327w(0) <= y_prenodeone_12_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9145w(0) <= y_prenodeone_12_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9148w(0) <= y_prenodeone_12_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9150w(0) <= y_prenodeone_12_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9152w(0) <= y_prenodeone_12_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9154w(0) <= y_prenodeone_12_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9156w(0) <= y_prenodeone_12_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9158w(0) <= y_prenodeone_12_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9210w(0) <= y_prenodeone_12_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9160w(0) <= y_prenodeone_12_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9162w(0) <= y_prenodeone_12_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9164w(0) <= y_prenodeone_12_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9166w(0) <= y_prenodeone_12_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9216w(0) <= y_prenodeone_12_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9222w(0) <= y_prenodeone_12_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9228w(0) <= y_prenodeone_12_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9234w(0) <= y_prenodeone_12_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9240w(0) <= y_prenodeone_12_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9246w(0) <= y_prenodeone_12_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range9252w(0) <= y_prenodeone_12_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10005w(0) <= y_prenodeone_13_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10064w(0) <= y_prenodeone_13_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10070w(0) <= y_prenodeone_13_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10076w(0) <= y_prenodeone_13_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10082w(0) <= y_prenodeone_13_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10088w(0) <= y_prenodeone_13_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10094w(0) <= y_prenodeone_13_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10100w(0) <= y_prenodeone_13_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10106w(0) <= y_prenodeone_13_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10112w(0) <= y_prenodeone_13_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10118w(0) <= y_prenodeone_13_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10010w(0) <= y_prenodeone_13_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10124w(0) <= y_prenodeone_13_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10127w(0) <= y_prenodeone_13_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9947w(0) <= y_prenodeone_13_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9950w(0) <= y_prenodeone_13_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9952w(0) <= y_prenodeone_13_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9954w(0) <= y_prenodeone_13_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9956w(0) <= y_prenodeone_13_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9958w(0) <= y_prenodeone_13_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9960w(0) <= y_prenodeone_13_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9962w(0) <= y_prenodeone_13_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10016w(0) <= y_prenodeone_13_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9964w(0) <= y_prenodeone_13_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9966w(0) <= y_prenodeone_13_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9968w(0) <= y_prenodeone_13_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9970w(0) <= y_prenodeone_13_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10022w(0) <= y_prenodeone_13_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10028w(0) <= y_prenodeone_13_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10034w(0) <= y_prenodeone_13_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10040w(0) <= y_prenodeone_13_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10046w(0) <= y_prenodeone_13_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10052w(0) <= y_prenodeone_13_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range10058w(0) <= y_prenodeone_13_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range864w(0) <= y_prenodeone_2_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range923w(0) <= y_prenodeone_2_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range929w(0) <= y_prenodeone_2_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range935w(0) <= y_prenodeone_2_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range941w(0) <= y_prenodeone_2_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range947w(0) <= y_prenodeone_2_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range953w(0) <= y_prenodeone_2_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range959w(0) <= y_prenodeone_2_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range965w(0) <= y_prenodeone_2_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range971w(0) <= y_prenodeone_2_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range977w(0) <= y_prenodeone_2_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range869w(0) <= y_prenodeone_2_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range983w(0) <= y_prenodeone_2_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range989w(0) <= y_prenodeone_2_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range995w(0) <= y_prenodeone_2_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1001w(0) <= y_prenodeone_2_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1007w(0) <= y_prenodeone_2_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1013w(0) <= y_prenodeone_2_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1019w(0) <= y_prenodeone_2_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1025w(0) <= y_prenodeone_2_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1031w(0) <= y_prenodeone_2_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1037w(0) <= y_prenodeone_2_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range875w(0) <= y_prenodeone_2_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1043w(0) <= y_prenodeone_2_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1049w(0) <= y_prenodeone_2_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range1052w(0) <= y_prenodeone_2_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range850w(0) <= y_prenodeone_2_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range881w(0) <= y_prenodeone_2_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range887w(0) <= y_prenodeone_2_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range893w(0) <= y_prenodeone_2_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range899w(0) <= y_prenodeone_2_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range905w(0) <= y_prenodeone_2_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range911w(0) <= y_prenodeone_2_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range917w(0) <= y_prenodeone_2_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1720w(0) <= y_prenodeone_3_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1779w(0) <= y_prenodeone_3_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1785w(0) <= y_prenodeone_3_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1791w(0) <= y_prenodeone_3_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1797w(0) <= y_prenodeone_3_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1803w(0) <= y_prenodeone_3_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1809w(0) <= y_prenodeone_3_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1815w(0) <= y_prenodeone_3_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1821w(0) <= y_prenodeone_3_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1827w(0) <= y_prenodeone_3_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1833w(0) <= y_prenodeone_3_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1725w(0) <= y_prenodeone_3_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1839w(0) <= y_prenodeone_3_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1845w(0) <= y_prenodeone_3_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1851w(0) <= y_prenodeone_3_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1857w(0) <= y_prenodeone_3_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1863w(0) <= y_prenodeone_3_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1869w(0) <= y_prenodeone_3_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1875w(0) <= y_prenodeone_3_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1881w(0) <= y_prenodeone_3_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1887w(0) <= y_prenodeone_3_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1893w(0) <= y_prenodeone_3_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1731w(0) <= y_prenodeone_3_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1899w(0) <= y_prenodeone_3_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1902w(0) <= y_prenodeone_3_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1702w(0) <= y_prenodeone_3_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1705w(0) <= y_prenodeone_3_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1737w(0) <= y_prenodeone_3_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1743w(0) <= y_prenodeone_3_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1749w(0) <= y_prenodeone_3_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1755w(0) <= y_prenodeone_3_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1761w(0) <= y_prenodeone_3_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1767w(0) <= y_prenodeone_3_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1773w(0) <= y_prenodeone_3_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2571w(0) <= y_prenodeone_4_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2630w(0) <= y_prenodeone_4_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2636w(0) <= y_prenodeone_4_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2642w(0) <= y_prenodeone_4_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2648w(0) <= y_prenodeone_4_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2654w(0) <= y_prenodeone_4_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2660w(0) <= y_prenodeone_4_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2666w(0) <= y_prenodeone_4_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2672w(0) <= y_prenodeone_4_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2678w(0) <= y_prenodeone_4_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2684w(0) <= y_prenodeone_4_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2576w(0) <= y_prenodeone_4_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2690w(0) <= y_prenodeone_4_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2696w(0) <= y_prenodeone_4_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2702w(0) <= y_prenodeone_4_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2708w(0) <= y_prenodeone_4_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2714w(0) <= y_prenodeone_4_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2720w(0) <= y_prenodeone_4_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2726w(0) <= y_prenodeone_4_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2732w(0) <= y_prenodeone_4_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2738w(0) <= y_prenodeone_4_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2744w(0) <= y_prenodeone_4_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2582w(0) <= y_prenodeone_4_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2747w(0) <= y_prenodeone_4_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2549w(0) <= y_prenodeone_4_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2552w(0) <= y_prenodeone_4_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2554w(0) <= y_prenodeone_4_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2588w(0) <= y_prenodeone_4_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2594w(0) <= y_prenodeone_4_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2600w(0) <= y_prenodeone_4_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2606w(0) <= y_prenodeone_4_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2612w(0) <= y_prenodeone_4_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2618w(0) <= y_prenodeone_4_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2624w(0) <= y_prenodeone_4_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3417w(0) <= y_prenodeone_5_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3476w(0) <= y_prenodeone_5_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3482w(0) <= y_prenodeone_5_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3488w(0) <= y_prenodeone_5_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3494w(0) <= y_prenodeone_5_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3500w(0) <= y_prenodeone_5_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3506w(0) <= y_prenodeone_5_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3512w(0) <= y_prenodeone_5_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3518w(0) <= y_prenodeone_5_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3524w(0) <= y_prenodeone_5_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3530w(0) <= y_prenodeone_5_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3422w(0) <= y_prenodeone_5_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3536w(0) <= y_prenodeone_5_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3542w(0) <= y_prenodeone_5_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3548w(0) <= y_prenodeone_5_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3554w(0) <= y_prenodeone_5_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3560w(0) <= y_prenodeone_5_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3566w(0) <= y_prenodeone_5_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3572w(0) <= y_prenodeone_5_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3578w(0) <= y_prenodeone_5_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3584w(0) <= y_prenodeone_5_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3587w(0) <= y_prenodeone_5_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3428w(0) <= y_prenodeone_5_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3391w(0) <= y_prenodeone_5_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3394w(0) <= y_prenodeone_5_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3396w(0) <= y_prenodeone_5_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3398w(0) <= y_prenodeone_5_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3434w(0) <= y_prenodeone_5_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3440w(0) <= y_prenodeone_5_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3446w(0) <= y_prenodeone_5_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3452w(0) <= y_prenodeone_5_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3458w(0) <= y_prenodeone_5_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3464w(0) <= y_prenodeone_5_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3470w(0) <= y_prenodeone_5_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4258w(0) <= y_prenodeone_6_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4317w(0) <= y_prenodeone_6_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4323w(0) <= y_prenodeone_6_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4329w(0) <= y_prenodeone_6_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4335w(0) <= y_prenodeone_6_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4341w(0) <= y_prenodeone_6_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4347w(0) <= y_prenodeone_6_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4353w(0) <= y_prenodeone_6_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4359w(0) <= y_prenodeone_6_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4365w(0) <= y_prenodeone_6_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4371w(0) <= y_prenodeone_6_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4263w(0) <= y_prenodeone_6_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4377w(0) <= y_prenodeone_6_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4383w(0) <= y_prenodeone_6_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4389w(0) <= y_prenodeone_6_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4395w(0) <= y_prenodeone_6_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4401w(0) <= y_prenodeone_6_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4407w(0) <= y_prenodeone_6_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4413w(0) <= y_prenodeone_6_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4419w(0) <= y_prenodeone_6_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4422w(0) <= y_prenodeone_6_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4228w(0) <= y_prenodeone_6_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4269w(0) <= y_prenodeone_6_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4231w(0) <= y_prenodeone_6_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4233w(0) <= y_prenodeone_6_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4235w(0) <= y_prenodeone_6_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4237w(0) <= y_prenodeone_6_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4275w(0) <= y_prenodeone_6_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4281w(0) <= y_prenodeone_6_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4287w(0) <= y_prenodeone_6_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4293w(0) <= y_prenodeone_6_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4299w(0) <= y_prenodeone_6_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4305w(0) <= y_prenodeone_6_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4311w(0) <= y_prenodeone_6_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5094w(0) <= y_prenodeone_7_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5153w(0) <= y_prenodeone_7_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5159w(0) <= y_prenodeone_7_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5165w(0) <= y_prenodeone_7_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5171w(0) <= y_prenodeone_7_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5177w(0) <= y_prenodeone_7_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5183w(0) <= y_prenodeone_7_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5189w(0) <= y_prenodeone_7_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5195w(0) <= y_prenodeone_7_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5201w(0) <= y_prenodeone_7_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5207w(0) <= y_prenodeone_7_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5099w(0) <= y_prenodeone_7_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5213w(0) <= y_prenodeone_7_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5219w(0) <= y_prenodeone_7_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5225w(0) <= y_prenodeone_7_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5231w(0) <= y_prenodeone_7_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5237w(0) <= y_prenodeone_7_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5243w(0) <= y_prenodeone_7_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5249w(0) <= y_prenodeone_7_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5252w(0) <= y_prenodeone_7_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5060w(0) <= y_prenodeone_7_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5063w(0) <= y_prenodeone_7_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5105w(0) <= y_prenodeone_7_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5065w(0) <= y_prenodeone_7_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5067w(0) <= y_prenodeone_7_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5069w(0) <= y_prenodeone_7_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5071w(0) <= y_prenodeone_7_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5111w(0) <= y_prenodeone_7_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5117w(0) <= y_prenodeone_7_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5123w(0) <= y_prenodeone_7_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5129w(0) <= y_prenodeone_7_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5135w(0) <= y_prenodeone_7_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5141w(0) <= y_prenodeone_7_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range5147w(0) <= y_prenodeone_7_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5925w(0) <= y_prenodeone_8_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5984w(0) <= y_prenodeone_8_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5990w(0) <= y_prenodeone_8_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5996w(0) <= y_prenodeone_8_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6002w(0) <= y_prenodeone_8_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6008w(0) <= y_prenodeone_8_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6014w(0) <= y_prenodeone_8_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6020w(0) <= y_prenodeone_8_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6026w(0) <= y_prenodeone_8_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6032w(0) <= y_prenodeone_8_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6038w(0) <= y_prenodeone_8_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5930w(0) <= y_prenodeone_8_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6044w(0) <= y_prenodeone_8_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6050w(0) <= y_prenodeone_8_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6056w(0) <= y_prenodeone_8_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6062w(0) <= y_prenodeone_8_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6068w(0) <= y_prenodeone_8_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6074w(0) <= y_prenodeone_8_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range6077w(0) <= y_prenodeone_8_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5887w(0) <= y_prenodeone_8_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5890w(0) <= y_prenodeone_8_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5892w(0) <= y_prenodeone_8_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5936w(0) <= y_prenodeone_8_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5894w(0) <= y_prenodeone_8_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5896w(0) <= y_prenodeone_8_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5898w(0) <= y_prenodeone_8_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5900w(0) <= y_prenodeone_8_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5942w(0) <= y_prenodeone_8_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5948w(0) <= y_prenodeone_8_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5954w(0) <= y_prenodeone_8_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5960w(0) <= y_prenodeone_8_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5966w(0) <= y_prenodeone_8_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5972w(0) <= y_prenodeone_8_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5978w(0) <= y_prenodeone_8_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6751w(0) <= y_prenodeone_9_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6810w(0) <= y_prenodeone_9_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6816w(0) <= y_prenodeone_9_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6822w(0) <= y_prenodeone_9_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6828w(0) <= y_prenodeone_9_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6834w(0) <= y_prenodeone_9_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6840w(0) <= y_prenodeone_9_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6846w(0) <= y_prenodeone_9_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6852w(0) <= y_prenodeone_9_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6858w(0) <= y_prenodeone_9_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6864w(0) <= y_prenodeone_9_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6756w(0) <= y_prenodeone_9_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6870w(0) <= y_prenodeone_9_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6876w(0) <= y_prenodeone_9_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6882w(0) <= y_prenodeone_9_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6888w(0) <= y_prenodeone_9_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6894w(0) <= y_prenodeone_9_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6897w(0) <= y_prenodeone_9_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6709w(0) <= y_prenodeone_9_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6712w(0) <= y_prenodeone_9_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6714w(0) <= y_prenodeone_9_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6716w(0) <= y_prenodeone_9_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6762w(0) <= y_prenodeone_9_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6718w(0) <= y_prenodeone_9_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6720w(0) <= y_prenodeone_9_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6722w(0) <= y_prenodeone_9_w(32);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6724w(0) <= y_prenodeone_9_w(33);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6768w(0) <= y_prenodeone_9_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6774w(0) <= y_prenodeone_9_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6780w(0) <= y_prenodeone_9_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6786w(0) <= y_prenodeone_9_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6792w(0) <= y_prenodeone_9_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6798w(0) <= y_prenodeone_9_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6804w(0) <= y_prenodeone_9_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7715w(0) <= y_prenodetwo_10_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7744w(0) <= y_prenodetwo_10_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7747w(0) <= y_prenodetwo_10_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7750w(0) <= y_prenodetwo_10_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7753w(0) <= y_prenodetwo_10_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7756w(0) <= y_prenodetwo_10_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7759w(0) <= y_prenodetwo_10_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7762w(0) <= y_prenodetwo_10_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7765w(0) <= y_prenodetwo_10_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7768w(0) <= y_prenodetwo_10_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7771w(0) <= y_prenodetwo_10_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7717w(0) <= y_prenodetwo_10_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7774w(0) <= y_prenodetwo_10_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7777w(0) <= y_prenodetwo_10_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7780w(0) <= y_prenodetwo_10_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7546w(0) <= y_prenodetwo_10_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7549w(0) <= y_prenodetwo_10_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7551w(0) <= y_prenodetwo_10_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7553w(0) <= y_prenodetwo_10_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7555w(0) <= y_prenodetwo_10_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7557w(0) <= y_prenodetwo_10_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7559w(0) <= y_prenodetwo_10_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7720w(0) <= y_prenodetwo_10_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7561w(0) <= y_prenodetwo_10_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7563w(0) <= y_prenodetwo_10_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7565w(0) <= y_prenodetwo_10_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7567w(0) <= y_prenodetwo_10_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7723w(0) <= y_prenodetwo_10_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7726w(0) <= y_prenodetwo_10_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7729w(0) <= y_prenodetwo_10_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7732w(0) <= y_prenodetwo_10_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7735w(0) <= y_prenodetwo_10_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7738w(0) <= y_prenodetwo_10_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7741w(0) <= y_prenodetwo_10_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8525w(0) <= y_prenodetwo_11_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8554w(0) <= y_prenodetwo_11_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8557w(0) <= y_prenodetwo_11_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8560w(0) <= y_prenodetwo_11_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8563w(0) <= y_prenodetwo_11_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8566w(0) <= y_prenodetwo_11_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8569w(0) <= y_prenodetwo_11_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8572w(0) <= y_prenodetwo_11_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8575w(0) <= y_prenodetwo_11_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8578w(0) <= y_prenodetwo_11_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8581w(0) <= y_prenodetwo_11_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8527w(0) <= y_prenodetwo_11_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8584w(0) <= y_prenodetwo_11_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8587w(0) <= y_prenodetwo_11_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8360w(0) <= y_prenodetwo_11_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8363w(0) <= y_prenodetwo_11_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8365w(0) <= y_prenodetwo_11_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8367w(0) <= y_prenodetwo_11_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8369w(0) <= y_prenodetwo_11_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8371w(0) <= y_prenodetwo_11_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8373w(0) <= y_prenodetwo_11_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8375w(0) <= y_prenodetwo_11_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8530w(0) <= y_prenodetwo_11_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8377w(0) <= y_prenodetwo_11_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8379w(0) <= y_prenodetwo_11_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8381w(0) <= y_prenodetwo_11_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8383w(0) <= y_prenodetwo_11_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8533w(0) <= y_prenodetwo_11_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8536w(0) <= y_prenodetwo_11_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8539w(0) <= y_prenodetwo_11_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8542w(0) <= y_prenodetwo_11_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8545w(0) <= y_prenodetwo_11_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8548w(0) <= y_prenodetwo_11_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range8551w(0) <= y_prenodetwo_11_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9330w(0) <= y_prenodetwo_12_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9359w(0) <= y_prenodetwo_12_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9362w(0) <= y_prenodetwo_12_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9365w(0) <= y_prenodetwo_12_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9368w(0) <= y_prenodetwo_12_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9371w(0) <= y_prenodetwo_12_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9374w(0) <= y_prenodetwo_12_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9377w(0) <= y_prenodetwo_12_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9380w(0) <= y_prenodetwo_12_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9383w(0) <= y_prenodetwo_12_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9386w(0) <= y_prenodetwo_12_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9332w(0) <= y_prenodetwo_12_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9389w(0) <= y_prenodetwo_12_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9169w(0) <= y_prenodetwo_12_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9172w(0) <= y_prenodetwo_12_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9174w(0) <= y_prenodetwo_12_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9176w(0) <= y_prenodetwo_12_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9178w(0) <= y_prenodetwo_12_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9180w(0) <= y_prenodetwo_12_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9182w(0) <= y_prenodetwo_12_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9184w(0) <= y_prenodetwo_12_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9186w(0) <= y_prenodetwo_12_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9335w(0) <= y_prenodetwo_12_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9188w(0) <= y_prenodetwo_12_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9190w(0) <= y_prenodetwo_12_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9192w(0) <= y_prenodetwo_12_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9194w(0) <= y_prenodetwo_12_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9338w(0) <= y_prenodetwo_12_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9341w(0) <= y_prenodetwo_12_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9344w(0) <= y_prenodetwo_12_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9347w(0) <= y_prenodetwo_12_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9350w(0) <= y_prenodetwo_12_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9353w(0) <= y_prenodetwo_12_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range9356w(0) <= y_prenodetwo_12_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10130w(0) <= y_prenodetwo_13_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10159w(0) <= y_prenodetwo_13_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10162w(0) <= y_prenodetwo_13_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10165w(0) <= y_prenodetwo_13_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10168w(0) <= y_prenodetwo_13_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10171w(0) <= y_prenodetwo_13_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10174w(0) <= y_prenodetwo_13_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10177w(0) <= y_prenodetwo_13_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10180w(0) <= y_prenodetwo_13_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10183w(0) <= y_prenodetwo_13_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10186w(0) <= y_prenodetwo_13_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10132w(0) <= y_prenodetwo_13_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9973w(0) <= y_prenodetwo_13_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9976w(0) <= y_prenodetwo_13_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9978w(0) <= y_prenodetwo_13_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9980w(0) <= y_prenodetwo_13_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9982w(0) <= y_prenodetwo_13_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9984w(0) <= y_prenodetwo_13_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9986w(0) <= y_prenodetwo_13_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9988w(0) <= y_prenodetwo_13_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9990w(0) <= y_prenodetwo_13_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9992w(0) <= y_prenodetwo_13_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10135w(0) <= y_prenodetwo_13_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9994w(0) <= y_prenodetwo_13_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9996w(0) <= y_prenodetwo_13_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9998w(0) <= y_prenodetwo_13_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10000w(0) <= y_prenodetwo_13_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10138w(0) <= y_prenodetwo_13_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10141w(0) <= y_prenodetwo_13_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10144w(0) <= y_prenodetwo_13_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10147w(0) <= y_prenodetwo_13_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10150w(0) <= y_prenodetwo_13_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10153w(0) <= y_prenodetwo_13_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range10156w(0) <= y_prenodetwo_13_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1055w(0) <= y_prenodetwo_2_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1084w(0) <= y_prenodetwo_2_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1087w(0) <= y_prenodetwo_2_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1090w(0) <= y_prenodetwo_2_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1093w(0) <= y_prenodetwo_2_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1096w(0) <= y_prenodetwo_2_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1099w(0) <= y_prenodetwo_2_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1102w(0) <= y_prenodetwo_2_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1105w(0) <= y_prenodetwo_2_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1108w(0) <= y_prenodetwo_2_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1111w(0) <= y_prenodetwo_2_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1057w(0) <= y_prenodetwo_2_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1114w(0) <= y_prenodetwo_2_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1117w(0) <= y_prenodetwo_2_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1120w(0) <= y_prenodetwo_2_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1123w(0) <= y_prenodetwo_2_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1126w(0) <= y_prenodetwo_2_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1129w(0) <= y_prenodetwo_2_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1132w(0) <= y_prenodetwo_2_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1135w(0) <= y_prenodetwo_2_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1138w(0) <= y_prenodetwo_2_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1141w(0) <= y_prenodetwo_2_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1060w(0) <= y_prenodetwo_2_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1144w(0) <= y_prenodetwo_2_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range854w(0) <= y_prenodetwo_2_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range857w(0) <= y_prenodetwo_2_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range859w(0) <= y_prenodetwo_2_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1063w(0) <= y_prenodetwo_2_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1066w(0) <= y_prenodetwo_2_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1069w(0) <= y_prenodetwo_2_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1072w(0) <= y_prenodetwo_2_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1075w(0) <= y_prenodetwo_2_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1078w(0) <= y_prenodetwo_2_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range1081w(0) <= y_prenodetwo_2_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1905w(0) <= y_prenodetwo_3_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1934w(0) <= y_prenodetwo_3_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1937w(0) <= y_prenodetwo_3_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1940w(0) <= y_prenodetwo_3_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1943w(0) <= y_prenodetwo_3_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1946w(0) <= y_prenodetwo_3_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1949w(0) <= y_prenodetwo_3_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1952w(0) <= y_prenodetwo_3_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1955w(0) <= y_prenodetwo_3_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1958w(0) <= y_prenodetwo_3_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1961w(0) <= y_prenodetwo_3_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1907w(0) <= y_prenodetwo_3_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1964w(0) <= y_prenodetwo_3_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1967w(0) <= y_prenodetwo_3_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1970w(0) <= y_prenodetwo_3_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1973w(0) <= y_prenodetwo_3_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1976w(0) <= y_prenodetwo_3_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1979w(0) <= y_prenodetwo_3_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1982w(0) <= y_prenodetwo_3_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1985w(0) <= y_prenodetwo_3_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1988w(0) <= y_prenodetwo_3_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1991w(0) <= y_prenodetwo_3_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1910w(0) <= y_prenodetwo_3_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1708w(0) <= y_prenodetwo_3_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1711w(0) <= y_prenodetwo_3_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1713w(0) <= y_prenodetwo_3_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1715w(0) <= y_prenodetwo_3_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1913w(0) <= y_prenodetwo_3_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1916w(0) <= y_prenodetwo_3_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1919w(0) <= y_prenodetwo_3_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1922w(0) <= y_prenodetwo_3_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1925w(0) <= y_prenodetwo_3_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1928w(0) <= y_prenodetwo_3_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1931w(0) <= y_prenodetwo_3_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2750w(0) <= y_prenodetwo_4_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2779w(0) <= y_prenodetwo_4_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2782w(0) <= y_prenodetwo_4_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2785w(0) <= y_prenodetwo_4_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2788w(0) <= y_prenodetwo_4_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2791w(0) <= y_prenodetwo_4_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2794w(0) <= y_prenodetwo_4_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2797w(0) <= y_prenodetwo_4_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2800w(0) <= y_prenodetwo_4_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2803w(0) <= y_prenodetwo_4_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2806w(0) <= y_prenodetwo_4_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2752w(0) <= y_prenodetwo_4_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2809w(0) <= y_prenodetwo_4_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2812w(0) <= y_prenodetwo_4_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2815w(0) <= y_prenodetwo_4_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2818w(0) <= y_prenodetwo_4_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2821w(0) <= y_prenodetwo_4_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2824w(0) <= y_prenodetwo_4_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2827w(0) <= y_prenodetwo_4_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2830w(0) <= y_prenodetwo_4_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2833w(0) <= y_prenodetwo_4_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2557w(0) <= y_prenodetwo_4_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2755w(0) <= y_prenodetwo_4_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2560w(0) <= y_prenodetwo_4_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2562w(0) <= y_prenodetwo_4_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2564w(0) <= y_prenodetwo_4_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2566w(0) <= y_prenodetwo_4_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2758w(0) <= y_prenodetwo_4_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2761w(0) <= y_prenodetwo_4_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2764w(0) <= y_prenodetwo_4_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2767w(0) <= y_prenodetwo_4_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2770w(0) <= y_prenodetwo_4_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2773w(0) <= y_prenodetwo_4_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2776w(0) <= y_prenodetwo_4_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3590w(0) <= y_prenodetwo_5_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3619w(0) <= y_prenodetwo_5_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3622w(0) <= y_prenodetwo_5_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3625w(0) <= y_prenodetwo_5_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3628w(0) <= y_prenodetwo_5_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3631w(0) <= y_prenodetwo_5_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3634w(0) <= y_prenodetwo_5_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3637w(0) <= y_prenodetwo_5_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3640w(0) <= y_prenodetwo_5_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3643w(0) <= y_prenodetwo_5_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3646w(0) <= y_prenodetwo_5_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3592w(0) <= y_prenodetwo_5_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3649w(0) <= y_prenodetwo_5_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3652w(0) <= y_prenodetwo_5_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3655w(0) <= y_prenodetwo_5_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3658w(0) <= y_prenodetwo_5_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3661w(0) <= y_prenodetwo_5_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3664w(0) <= y_prenodetwo_5_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3667w(0) <= y_prenodetwo_5_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3670w(0) <= y_prenodetwo_5_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3401w(0) <= y_prenodetwo_5_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3404w(0) <= y_prenodetwo_5_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3595w(0) <= y_prenodetwo_5_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3406w(0) <= y_prenodetwo_5_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3408w(0) <= y_prenodetwo_5_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3410w(0) <= y_prenodetwo_5_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3412w(0) <= y_prenodetwo_5_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3598w(0) <= y_prenodetwo_5_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3601w(0) <= y_prenodetwo_5_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3604w(0) <= y_prenodetwo_5_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3607w(0) <= y_prenodetwo_5_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3610w(0) <= y_prenodetwo_5_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3613w(0) <= y_prenodetwo_5_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3616w(0) <= y_prenodetwo_5_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4425w(0) <= y_prenodetwo_6_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4454w(0) <= y_prenodetwo_6_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4457w(0) <= y_prenodetwo_6_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4460w(0) <= y_prenodetwo_6_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4463w(0) <= y_prenodetwo_6_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4466w(0) <= y_prenodetwo_6_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4469w(0) <= y_prenodetwo_6_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4472w(0) <= y_prenodetwo_6_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4475w(0) <= y_prenodetwo_6_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4478w(0) <= y_prenodetwo_6_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4481w(0) <= y_prenodetwo_6_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4427w(0) <= y_prenodetwo_6_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4484w(0) <= y_prenodetwo_6_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4487w(0) <= y_prenodetwo_6_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4490w(0) <= y_prenodetwo_6_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4493w(0) <= y_prenodetwo_6_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4496w(0) <= y_prenodetwo_6_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4499w(0) <= y_prenodetwo_6_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4502w(0) <= y_prenodetwo_6_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4240w(0) <= y_prenodetwo_6_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4243w(0) <= y_prenodetwo_6_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4245w(0) <= y_prenodetwo_6_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4430w(0) <= y_prenodetwo_6_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4247w(0) <= y_prenodetwo_6_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4249w(0) <= y_prenodetwo_6_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4251w(0) <= y_prenodetwo_6_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4253w(0) <= y_prenodetwo_6_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4433w(0) <= y_prenodetwo_6_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4436w(0) <= y_prenodetwo_6_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4439w(0) <= y_prenodetwo_6_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4442w(0) <= y_prenodetwo_6_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4445w(0) <= y_prenodetwo_6_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4448w(0) <= y_prenodetwo_6_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4451w(0) <= y_prenodetwo_6_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5255w(0) <= y_prenodetwo_7_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5284w(0) <= y_prenodetwo_7_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5287w(0) <= y_prenodetwo_7_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5290w(0) <= y_prenodetwo_7_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5293w(0) <= y_prenodetwo_7_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5296w(0) <= y_prenodetwo_7_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5299w(0) <= y_prenodetwo_7_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5302w(0) <= y_prenodetwo_7_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5305w(0) <= y_prenodetwo_7_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5308w(0) <= y_prenodetwo_7_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5311w(0) <= y_prenodetwo_7_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5257w(0) <= y_prenodetwo_7_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5314w(0) <= y_prenodetwo_7_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5317w(0) <= y_prenodetwo_7_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5320w(0) <= y_prenodetwo_7_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5323w(0) <= y_prenodetwo_7_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5326w(0) <= y_prenodetwo_7_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5329w(0) <= y_prenodetwo_7_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5074w(0) <= y_prenodetwo_7_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5077w(0) <= y_prenodetwo_7_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5079w(0) <= y_prenodetwo_7_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5081w(0) <= y_prenodetwo_7_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5260w(0) <= y_prenodetwo_7_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5083w(0) <= y_prenodetwo_7_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5085w(0) <= y_prenodetwo_7_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5087w(0) <= y_prenodetwo_7_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5089w(0) <= y_prenodetwo_7_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5263w(0) <= y_prenodetwo_7_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5266w(0) <= y_prenodetwo_7_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5269w(0) <= y_prenodetwo_7_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5272w(0) <= y_prenodetwo_7_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5275w(0) <= y_prenodetwo_7_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5278w(0) <= y_prenodetwo_7_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range5281w(0) <= y_prenodetwo_7_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6080w(0) <= y_prenodetwo_8_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6109w(0) <= y_prenodetwo_8_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6112w(0) <= y_prenodetwo_8_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6115w(0) <= y_prenodetwo_8_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6118w(0) <= y_prenodetwo_8_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6121w(0) <= y_prenodetwo_8_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6124w(0) <= y_prenodetwo_8_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6127w(0) <= y_prenodetwo_8_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6130w(0) <= y_prenodetwo_8_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6133w(0) <= y_prenodetwo_8_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6136w(0) <= y_prenodetwo_8_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6082w(0) <= y_prenodetwo_8_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6139w(0) <= y_prenodetwo_8_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6142w(0) <= y_prenodetwo_8_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6145w(0) <= y_prenodetwo_8_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6148w(0) <= y_prenodetwo_8_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6151w(0) <= y_prenodetwo_8_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5903w(0) <= y_prenodetwo_8_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5906w(0) <= y_prenodetwo_8_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5908w(0) <= y_prenodetwo_8_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5910w(0) <= y_prenodetwo_8_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5912w(0) <= y_prenodetwo_8_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6085w(0) <= y_prenodetwo_8_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5914w(0) <= y_prenodetwo_8_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5916w(0) <= y_prenodetwo_8_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5918w(0) <= y_prenodetwo_8_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5920w(0) <= y_prenodetwo_8_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6088w(0) <= y_prenodetwo_8_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6091w(0) <= y_prenodetwo_8_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6094w(0) <= y_prenodetwo_8_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6097w(0) <= y_prenodetwo_8_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6100w(0) <= y_prenodetwo_8_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6103w(0) <= y_prenodetwo_8_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range6106w(0) <= y_prenodetwo_8_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6900w(0) <= y_prenodetwo_9_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6929w(0) <= y_prenodetwo_9_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6932w(0) <= y_prenodetwo_9_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6935w(0) <= y_prenodetwo_9_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6938w(0) <= y_prenodetwo_9_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6941w(0) <= y_prenodetwo_9_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6944w(0) <= y_prenodetwo_9_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6947w(0) <= y_prenodetwo_9_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6950w(0) <= y_prenodetwo_9_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6953w(0) <= y_prenodetwo_9_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6956w(0) <= y_prenodetwo_9_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6902w(0) <= y_prenodetwo_9_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6959w(0) <= y_prenodetwo_9_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6962w(0) <= y_prenodetwo_9_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6965w(0) <= y_prenodetwo_9_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6968w(0) <= y_prenodetwo_9_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6727w(0) <= y_prenodetwo_9_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6730w(0) <= y_prenodetwo_9_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6732w(0) <= y_prenodetwo_9_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6734w(0) <= y_prenodetwo_9_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6736w(0) <= y_prenodetwo_9_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6738w(0) <= y_prenodetwo_9_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6905w(0) <= y_prenodetwo_9_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6740w(0) <= y_prenodetwo_9_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6742w(0) <= y_prenodetwo_9_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6744w(0) <= y_prenodetwo_9_w(32);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6746w(0) <= y_prenodetwo_9_w(33);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6908w(0) <= y_prenodetwo_9_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6911w(0) <= y_prenodetwo_9_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6914w(0) <= y_prenodetwo_9_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6917w(0) <= y_prenodetwo_9_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6920w(0) <= y_prenodetwo_9_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6923w(0) <= y_prenodetwo_9_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6926w(0) <= y_prenodetwo_9_w(9);
	cata_0_cordic_atan :  sinhw_altfp_sincos_cordic_atan_45b
	  PORT MAP ( 
		arctan => wire_cata_0_cordic_atan_arctan,
		indexbit => indexbitff(0)
	  );
	cata_10_cordic_atan :  sinhw_altfp_sincos_cordic_atan_l6b
	  PORT MAP ( 
		arctan => wire_cata_10_cordic_atan_arctan,
		indexbit => indexbitff(10)
	  );
	cata_11_cordic_atan :  sinhw_altfp_sincos_cordic_atan_m6b
	  PORT MAP ( 
		arctan => wire_cata_11_cordic_atan_arctan,
		indexbit => indexbitff(11)
	  );
	cata_12_cordic_atan :  sinhw_altfp_sincos_cordic_atan_n6b
	  PORT MAP ( 
		arctan => wire_cata_12_cordic_atan_arctan,
		indexbit => indexbitff(12)
	  );
	cata_13_cordic_atan :  sinhw_altfp_sincos_cordic_atan_o6b
	  PORT MAP ( 
		arctan => wire_cata_13_cordic_atan_arctan,
		indexbit => indexbitff(13)
	  );
	cata_1_cordic_atan :  sinhw_altfp_sincos_cordic_atan_55b
	  PORT MAP ( 
		arctan => wire_cata_1_cordic_atan_arctan,
		indexbit => indexbitff(1)
	  );
	cata_2_cordic_atan :  sinhw_altfp_sincos_cordic_atan_65b
	  PORT MAP ( 
		arctan => wire_cata_2_cordic_atan_arctan,
		indexbit => indexbitff(2)
	  );
	cata_3_cordic_atan :  sinhw_altfp_sincos_cordic_atan_75b
	  PORT MAP ( 
		arctan => wire_cata_3_cordic_atan_arctan,
		indexbit => indexbitff(3)
	  );
	cata_4_cordic_atan :  sinhw_altfp_sincos_cordic_atan_85b
	  PORT MAP ( 
		arctan => wire_cata_4_cordic_atan_arctan,
		indexbit => indexbitff(4)
	  );
	cata_5_cordic_atan :  sinhw_altfp_sincos_cordic_atan_95b
	  PORT MAP ( 
		arctan => wire_cata_5_cordic_atan_arctan,
		indexbit => indexbitff(5)
	  );
	cata_6_cordic_atan :  sinhw_altfp_sincos_cordic_atan_a5b
	  PORT MAP ( 
		arctan => wire_cata_6_cordic_atan_arctan,
		indexbit => indexbitff(6)
	  );
	cata_7_cordic_atan :  sinhw_altfp_sincos_cordic_atan_b5b
	  PORT MAP ( 
		arctan => wire_cata_7_cordic_atan_arctan,
		indexbit => indexbitff(7)
	  );
	cata_8_cordic_atan :  sinhw_altfp_sincos_cordic_atan_c5b
	  PORT MAP ( 
		arctan => wire_cata_8_cordic_atan_arctan,
		indexbit => indexbitff(8)
	  );
	cata_9_cordic_atan :  sinhw_altfp_sincos_cordic_atan_d5b
	  PORT MAP ( 
		arctan => wire_cata_9_cordic_atan_arctan,
		indexbit => indexbitff(9)
	  );
	cxs :  sinhw_altfp_sincos_cordic_start_709
	  PORT MAP ( 
		index => startindex_w,
		value => wire_cxs_value
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cdaff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cdaff_0 <= delay_input_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cdaff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cdaff_1 <= cdaff_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cdaff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cdaff_2 <= cdaff_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN indexbitff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN indexbitff <= ( indexbitff(15 DOWNTO 0) & indexbit);
			END IF;
		END IF;
	END PROCESS;
	wire_indexbitff_w_lg_w_q_range581w679w(0) <= NOT wire_indexbitff_w_q_range581w(0);
	wire_indexbitff_w_lg_w_q_range610w8590w(0) <= NOT wire_indexbitff_w_q_range610w(0);
	wire_indexbitff_w_lg_w_q_range613w9392w(0) <= NOT wire_indexbitff_w_q_range613w(0);
	wire_indexbitff_w_lg_w_q_range616w10189w(0) <= NOT wire_indexbitff_w_q_range616w(0);
	wire_indexbitff_w_lg_w_q_range10749w10752w(0) <= NOT wire_indexbitff_w_q_range10749w(0);
	wire_indexbitff_w_lg_w_q_range583w1147w(0) <= NOT wire_indexbitff_w_q_range583w(0);
	wire_indexbitff_w_lg_w_q_range586w1994w(0) <= NOT wire_indexbitff_w_q_range586w(0);
	wire_indexbitff_w_lg_w_q_range589w2836w(0) <= NOT wire_indexbitff_w_q_range589w(0);
	wire_indexbitff_w_lg_w_q_range592w3673w(0) <= NOT wire_indexbitff_w_q_range592w(0);
	wire_indexbitff_w_lg_w_q_range595w4505w(0) <= NOT wire_indexbitff_w_q_range595w(0);
	wire_indexbitff_w_lg_w_q_range598w5332w(0) <= NOT wire_indexbitff_w_q_range598w(0);
	wire_indexbitff_w_lg_w_q_range601w6154w(0) <= NOT wire_indexbitff_w_q_range601w(0);
	wire_indexbitff_w_lg_w_q_range604w6971w(0) <= NOT wire_indexbitff_w_q_range604w(0);
	wire_indexbitff_w_lg_w_q_range607w7783w(0) <= NOT wire_indexbitff_w_q_range607w(0);
	wire_indexbitff_w_q_range581w(0) <= indexbitff(0);
	wire_indexbitff_w_q_range610w(0) <= indexbitff(10);
	wire_indexbitff_w_q_range613w(0) <= indexbitff(11);
	wire_indexbitff_w_q_range616w(0) <= indexbitff(12);
	wire_indexbitff_w_q_range10749w(0) <= indexbitff(16);
	wire_indexbitff_w_q_range583w(0) <= indexbitff(1);
	wire_indexbitff_w_q_range586w(0) <= indexbitff(2);
	wire_indexbitff_w_q_range589w(0) <= indexbitff(3);
	wire_indexbitff_w_q_range592w(0) <= indexbitff(4);
	wire_indexbitff_w_q_range595w(0) <= indexbitff(5);
	wire_indexbitff_w_q_range598w(0) <= indexbitff(6);
	wire_indexbitff_w_q_range601w(0) <= indexbitff(7);
	wire_indexbitff_w_q_range604w(0) <= indexbitff(8);
	wire_indexbitff_w_q_range607w(0) <= indexbitff(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sincosbitff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN sincosbitff <= ( sincosbitff(15 DOWNTO 0) & sincosbit);
			END IF;
		END IF;
	END PROCESS;
	wire_sincosbitff_w_lg_w_q_range668w10739w(0) <= NOT wire_sincosbitff_w_q_range668w(0);
	wire_sincosbitff_w_lg_w_q_range10746w10747w(0) <= NOT wire_sincosbitff_w_q_range10746w(0);
	wire_sincosbitff_w_q_range668w(0) <= sincosbitff(13);
	wire_sincosbitff_w_q_range10746w(0) <= sincosbitff(16);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sincosff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN sincosff <= wire_sincos_add_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_0 <= x_start_node_w;
			END IF;
		END IF;
	END PROCESS;
	wire_x_pipeff_0_w_lg_w_q_range680w681w(0) <= wire_x_pipeff_0_w_q_range680w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range721w733w(0) <= wire_x_pipeff_0_w_q_range721w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range721w722w(0) <= wire_x_pipeff_0_w_q_range721w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range726w738w(0) <= wire_x_pipeff_0_w_q_range726w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range726w727w(0) <= wire_x_pipeff_0_w_q_range726w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range731w743w(0) <= wire_x_pipeff_0_w_q_range731w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range731w732w(0) <= wire_x_pipeff_0_w_q_range731w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range736w748w(0) <= wire_x_pipeff_0_w_q_range736w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range736w737w(0) <= wire_x_pipeff_0_w_q_range736w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range741w753w(0) <= wire_x_pipeff_0_w_q_range741w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range741w742w(0) <= wire_x_pipeff_0_w_q_range741w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range746w758w(0) <= wire_x_pipeff_0_w_q_range746w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range746w747w(0) <= wire_x_pipeff_0_w_q_range746w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range751w763w(0) <= wire_x_pipeff_0_w_q_range751w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range751w752w(0) <= wire_x_pipeff_0_w_q_range751w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range756w768w(0) <= wire_x_pipeff_0_w_q_range756w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range756w757w(0) <= wire_x_pipeff_0_w_q_range756w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range761w773w(0) <= wire_x_pipeff_0_w_q_range761w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range761w762w(0) <= wire_x_pipeff_0_w_q_range761w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range766w778w(0) <= wire_x_pipeff_0_w_q_range766w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range766w767w(0) <= wire_x_pipeff_0_w_q_range766w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range687w688w(0) <= wire_x_pipeff_0_w_q_range687w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range771w783w(0) <= wire_x_pipeff_0_w_q_range771w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range771w772w(0) <= wire_x_pipeff_0_w_q_range771w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range776w788w(0) <= wire_x_pipeff_0_w_q_range776w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range776w777w(0) <= wire_x_pipeff_0_w_q_range776w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range781w793w(0) <= wire_x_pipeff_0_w_q_range781w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range781w782w(0) <= wire_x_pipeff_0_w_q_range781w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range786w798w(0) <= wire_x_pipeff_0_w_q_range786w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range786w787w(0) <= wire_x_pipeff_0_w_q_range786w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range791w803w(0) <= wire_x_pipeff_0_w_q_range791w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range791w792w(0) <= wire_x_pipeff_0_w_q_range791w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range796w808w(0) <= wire_x_pipeff_0_w_q_range796w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range796w797w(0) <= wire_x_pipeff_0_w_q_range796w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range801w813w(0) <= wire_x_pipeff_0_w_q_range801w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range801w802w(0) <= wire_x_pipeff_0_w_q_range801w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range806w818w(0) <= wire_x_pipeff_0_w_q_range806w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range806w807w(0) <= wire_x_pipeff_0_w_q_range806w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range811w823w(0) <= wire_x_pipeff_0_w_q_range811w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range811w812w(0) <= wire_x_pipeff_0_w_q_range811w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range816w828w(0) <= wire_x_pipeff_0_w_q_range816w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range816w817w(0) <= wire_x_pipeff_0_w_q_range816w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range677w693w(0) <= wire_x_pipeff_0_w_q_range677w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range677w678w(0) <= wire_x_pipeff_0_w_q_range677w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range821w833w(0) <= wire_x_pipeff_0_w_q_range821w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range821w822w(0) <= wire_x_pipeff_0_w_q_range821w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range826w838w(0) <= wire_x_pipeff_0_w_q_range826w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range826w827w(0) <= wire_x_pipeff_0_w_q_range826w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range831w841w(0) <= wire_x_pipeff_0_w_q_range831w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range831w832w(0) <= wire_x_pipeff_0_w_q_range831w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range836w837w(0) <= wire_x_pipeff_0_w_q_range836w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range685w698w(0) <= wire_x_pipeff_0_w_q_range685w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range685w686w(0) <= wire_x_pipeff_0_w_q_range685w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range691w703w(0) <= wire_x_pipeff_0_w_q_range691w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range691w692w(0) <= wire_x_pipeff_0_w_q_range691w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range696w708w(0) <= wire_x_pipeff_0_w_q_range696w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range696w697w(0) <= wire_x_pipeff_0_w_q_range696w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range701w713w(0) <= wire_x_pipeff_0_w_q_range701w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range701w702w(0) <= wire_x_pipeff_0_w_q_range701w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range706w718w(0) <= wire_x_pipeff_0_w_q_range706w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range706w707w(0) <= wire_x_pipeff_0_w_q_range706w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range711w723w(0) <= wire_x_pipeff_0_w_q_range711w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range711w712w(0) <= wire_x_pipeff_0_w_q_range711w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range716w728w(0) <= wire_x_pipeff_0_w_q_range716w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_q_range716w717w(0) <= wire_x_pipeff_0_w_q_range716w(0) AND wire_indexbitff_w_q_range581w(0);
	wire_x_pipeff_0_w_lg_w_q_range836w843w(0) <= wire_x_pipeff_0_w_q_range836w(0) AND wire_indexbitff_w_lg_w_q_range581w679w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range680w681w682w(0) <= wire_x_pipeff_0_w_lg_w_q_range680w681w(0) OR wire_x_pipeff_0_w_lg_w_q_range677w678w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range721w733w734w(0) <= wire_x_pipeff_0_w_lg_w_q_range721w733w(0) OR wire_x_pipeff_0_w_lg_w_q_range731w732w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range726w738w739w(0) <= wire_x_pipeff_0_w_lg_w_q_range726w738w(0) OR wire_x_pipeff_0_w_lg_w_q_range736w737w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range731w743w744w(0) <= wire_x_pipeff_0_w_lg_w_q_range731w743w(0) OR wire_x_pipeff_0_w_lg_w_q_range741w742w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range736w748w749w(0) <= wire_x_pipeff_0_w_lg_w_q_range736w748w(0) OR wire_x_pipeff_0_w_lg_w_q_range746w747w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range741w753w754w(0) <= wire_x_pipeff_0_w_lg_w_q_range741w753w(0) OR wire_x_pipeff_0_w_lg_w_q_range751w752w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range746w758w759w(0) <= wire_x_pipeff_0_w_lg_w_q_range746w758w(0) OR wire_x_pipeff_0_w_lg_w_q_range756w757w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range751w763w764w(0) <= wire_x_pipeff_0_w_lg_w_q_range751w763w(0) OR wire_x_pipeff_0_w_lg_w_q_range761w762w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range756w768w769w(0) <= wire_x_pipeff_0_w_lg_w_q_range756w768w(0) OR wire_x_pipeff_0_w_lg_w_q_range766w767w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range761w773w774w(0) <= wire_x_pipeff_0_w_lg_w_q_range761w773w(0) OR wire_x_pipeff_0_w_lg_w_q_range771w772w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range766w778w779w(0) <= wire_x_pipeff_0_w_lg_w_q_range766w778w(0) OR wire_x_pipeff_0_w_lg_w_q_range776w777w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range687w688w689w(0) <= wire_x_pipeff_0_w_lg_w_q_range687w688w(0) OR wire_x_pipeff_0_w_lg_w_q_range685w686w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range771w783w784w(0) <= wire_x_pipeff_0_w_lg_w_q_range771w783w(0) OR wire_x_pipeff_0_w_lg_w_q_range781w782w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range776w788w789w(0) <= wire_x_pipeff_0_w_lg_w_q_range776w788w(0) OR wire_x_pipeff_0_w_lg_w_q_range786w787w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range781w793w794w(0) <= wire_x_pipeff_0_w_lg_w_q_range781w793w(0) OR wire_x_pipeff_0_w_lg_w_q_range791w792w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range786w798w799w(0) <= wire_x_pipeff_0_w_lg_w_q_range786w798w(0) OR wire_x_pipeff_0_w_lg_w_q_range796w797w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range791w803w804w(0) <= wire_x_pipeff_0_w_lg_w_q_range791w803w(0) OR wire_x_pipeff_0_w_lg_w_q_range801w802w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range796w808w809w(0) <= wire_x_pipeff_0_w_lg_w_q_range796w808w(0) OR wire_x_pipeff_0_w_lg_w_q_range806w807w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range801w813w814w(0) <= wire_x_pipeff_0_w_lg_w_q_range801w813w(0) OR wire_x_pipeff_0_w_lg_w_q_range811w812w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range806w818w819w(0) <= wire_x_pipeff_0_w_lg_w_q_range806w818w(0) OR wire_x_pipeff_0_w_lg_w_q_range816w817w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range811w823w824w(0) <= wire_x_pipeff_0_w_lg_w_q_range811w823w(0) OR wire_x_pipeff_0_w_lg_w_q_range821w822w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range816w828w829w(0) <= wire_x_pipeff_0_w_lg_w_q_range816w828w(0) OR wire_x_pipeff_0_w_lg_w_q_range826w827w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range677w693w694w(0) <= wire_x_pipeff_0_w_lg_w_q_range677w693w(0) OR wire_x_pipeff_0_w_lg_w_q_range691w692w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range821w833w834w(0) <= wire_x_pipeff_0_w_lg_w_q_range821w833w(0) OR wire_x_pipeff_0_w_lg_w_q_range831w832w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range826w838w839w(0) <= wire_x_pipeff_0_w_lg_w_q_range826w838w(0) OR wire_x_pipeff_0_w_lg_w_q_range836w837w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range685w698w699w(0) <= wire_x_pipeff_0_w_lg_w_q_range685w698w(0) OR wire_x_pipeff_0_w_lg_w_q_range696w697w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range691w703w704w(0) <= wire_x_pipeff_0_w_lg_w_q_range691w703w(0) OR wire_x_pipeff_0_w_lg_w_q_range701w702w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range696w708w709w(0) <= wire_x_pipeff_0_w_lg_w_q_range696w708w(0) OR wire_x_pipeff_0_w_lg_w_q_range706w707w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range701w713w714w(0) <= wire_x_pipeff_0_w_lg_w_q_range701w713w(0) OR wire_x_pipeff_0_w_lg_w_q_range711w712w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range706w718w719w(0) <= wire_x_pipeff_0_w_lg_w_q_range706w718w(0) OR wire_x_pipeff_0_w_lg_w_q_range716w717w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range711w723w724w(0) <= wire_x_pipeff_0_w_lg_w_q_range711w723w(0) OR wire_x_pipeff_0_w_lg_w_q_range721w722w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range716w728w729w(0) <= wire_x_pipeff_0_w_lg_w_q_range716w728w(0) OR wire_x_pipeff_0_w_lg_w_q_range726w727w(0);
	wire_x_pipeff_0_w_q_range680w(0) <= x_pipeff_0(0);
	wire_x_pipeff_0_w_q_range721w(0) <= x_pipeff_0(10);
	wire_x_pipeff_0_w_q_range726w(0) <= x_pipeff_0(11);
	wire_x_pipeff_0_w_q_range731w(0) <= x_pipeff_0(12);
	wire_x_pipeff_0_w_q_range736w(0) <= x_pipeff_0(13);
	wire_x_pipeff_0_w_q_range741w(0) <= x_pipeff_0(14);
	wire_x_pipeff_0_w_q_range746w(0) <= x_pipeff_0(15);
	wire_x_pipeff_0_w_q_range751w(0) <= x_pipeff_0(16);
	wire_x_pipeff_0_w_q_range756w(0) <= x_pipeff_0(17);
	wire_x_pipeff_0_w_q_range761w(0) <= x_pipeff_0(18);
	wire_x_pipeff_0_w_q_range766w(0) <= x_pipeff_0(19);
	wire_x_pipeff_0_w_q_range687w(0) <= x_pipeff_0(1);
	wire_x_pipeff_0_w_q_range771w(0) <= x_pipeff_0(20);
	wire_x_pipeff_0_w_q_range776w(0) <= x_pipeff_0(21);
	wire_x_pipeff_0_w_q_range781w(0) <= x_pipeff_0(22);
	wire_x_pipeff_0_w_q_range786w(0) <= x_pipeff_0(23);
	wire_x_pipeff_0_w_q_range791w(0) <= x_pipeff_0(24);
	wire_x_pipeff_0_w_q_range796w(0) <= x_pipeff_0(25);
	wire_x_pipeff_0_w_q_range801w(0) <= x_pipeff_0(26);
	wire_x_pipeff_0_w_q_range806w(0) <= x_pipeff_0(27);
	wire_x_pipeff_0_w_q_range811w(0) <= x_pipeff_0(28);
	wire_x_pipeff_0_w_q_range816w(0) <= x_pipeff_0(29);
	wire_x_pipeff_0_w_q_range677w(0) <= x_pipeff_0(2);
	wire_x_pipeff_0_w_q_range821w(0) <= x_pipeff_0(30);
	wire_x_pipeff_0_w_q_range826w(0) <= x_pipeff_0(31);
	wire_x_pipeff_0_w_q_range831w(0) <= x_pipeff_0(32);
	wire_x_pipeff_0_w_q_range836w(0) <= x_pipeff_0(33);
	wire_x_pipeff_0_w_q_range685w(0) <= x_pipeff_0(3);
	wire_x_pipeff_0_w_q_range691w(0) <= x_pipeff_0(4);
	wire_x_pipeff_0_w_q_range696w(0) <= x_pipeff_0(5);
	wire_x_pipeff_0_w_q_range701w(0) <= x_pipeff_0(6);
	wire_x_pipeff_0_w_q_range706w(0) <= x_pipeff_0(7);
	wire_x_pipeff_0_w_q_range711w(0) <= x_pipeff_0(8);
	wire_x_pipeff_0_w_q_range716w(0) <= x_pipeff_0(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_1 <= x_pipeff_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_10 <= x_pipenode_10_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_11 <= x_pipenode_11_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_12 <= x_pipenode_12_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_13 <= x_pipenode_13_w;
			END IF;
		END IF;
	END PROCESS;
	loop32 : FOR i IN 0 TO 33 GENERATE 
		wire_x_pipeff_13_w_lg_q10744w(i) <= x_pipeff_13(i) AND wire_sincosbitff_w_lg_w_q_range668w10739w(0);
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 33 GENERATE 
		wire_x_pipeff_13_w_lg_q10741w(i) <= x_pipeff_13(i) AND wire_sincosbitff_w_q_range668w(0);
	END GENERATE loop33;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_2 <= x_pipenode_2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_3 <= x_pipenode_3_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_4 <= x_pipenode_4_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_5 <= x_pipenode_5_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_6 <= x_pipenode_6_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_7 <= x_pipenode_7_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_8 <= x_pipenode_8_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_9 <= x_pipenode_9_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(0) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(0) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(1) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(1) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(2) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(2) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(3) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(3) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(4) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(4) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(5) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(5) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(6) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(6) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(7) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(7) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(8) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(8) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(9) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(9) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(10) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(10) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(11) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(11) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(12) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(12) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(13) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(13) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(14) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(14) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(15) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(15) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(16) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(16) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(17) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(17) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(18) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(18) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(19) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(19) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(20) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(20) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(21) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(21) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(22) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(22) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(23) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(23) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(24) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(24) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(25) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(25) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(26) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(26) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(27) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(27) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(28) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(28) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(29) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(29) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(30) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(30) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(31) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(31) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(32) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(32) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(33) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(33) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_1 <= wire_y_pipeff1_add_result;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_1_w_lg_w_q_range913w914w(0) <= NOT wire_y_pipeff_1_w_q_range913w(0);
	wire_y_pipeff_1_w_lg_w_q_range919w920w(0) <= NOT wire_y_pipeff_1_w_q_range919w(0);
	wire_y_pipeff_1_w_lg_w_q_range925w926w(0) <= NOT wire_y_pipeff_1_w_q_range925w(0);
	wire_y_pipeff_1_w_lg_w_q_range931w932w(0) <= NOT wire_y_pipeff_1_w_q_range931w(0);
	wire_y_pipeff_1_w_lg_w_q_range937w938w(0) <= NOT wire_y_pipeff_1_w_q_range937w(0);
	wire_y_pipeff_1_w_lg_w_q_range943w944w(0) <= NOT wire_y_pipeff_1_w_q_range943w(0);
	wire_y_pipeff_1_w_lg_w_q_range949w950w(0) <= NOT wire_y_pipeff_1_w_q_range949w(0);
	wire_y_pipeff_1_w_lg_w_q_range955w956w(0) <= NOT wire_y_pipeff_1_w_q_range955w(0);
	wire_y_pipeff_1_w_lg_w_q_range961w962w(0) <= NOT wire_y_pipeff_1_w_q_range961w(0);
	wire_y_pipeff_1_w_lg_w_q_range967w968w(0) <= NOT wire_y_pipeff_1_w_q_range967w(0);
	wire_y_pipeff_1_w_lg_w_q_range860w861w(0) <= NOT wire_y_pipeff_1_w_q_range860w(0);
	wire_y_pipeff_1_w_lg_w_q_range973w974w(0) <= NOT wire_y_pipeff_1_w_q_range973w(0);
	wire_y_pipeff_1_w_lg_w_q_range979w980w(0) <= NOT wire_y_pipeff_1_w_q_range979w(0);
	wire_y_pipeff_1_w_lg_w_q_range985w986w(0) <= NOT wire_y_pipeff_1_w_q_range985w(0);
	wire_y_pipeff_1_w_lg_w_q_range991w992w(0) <= NOT wire_y_pipeff_1_w_q_range991w(0);
	wire_y_pipeff_1_w_lg_w_q_range997w998w(0) <= NOT wire_y_pipeff_1_w_q_range997w(0);
	wire_y_pipeff_1_w_lg_w_q_range1003w1004w(0) <= NOT wire_y_pipeff_1_w_q_range1003w(0);
	wire_y_pipeff_1_w_lg_w_q_range1009w1010w(0) <= NOT wire_y_pipeff_1_w_q_range1009w(0);
	wire_y_pipeff_1_w_lg_w_q_range1015w1016w(0) <= NOT wire_y_pipeff_1_w_q_range1015w(0);
	wire_y_pipeff_1_w_lg_w_q_range1021w1022w(0) <= NOT wire_y_pipeff_1_w_q_range1021w(0);
	wire_y_pipeff_1_w_lg_w_q_range1027w1028w(0) <= NOT wire_y_pipeff_1_w_q_range1027w(0);
	wire_y_pipeff_1_w_lg_w_q_range865w866w(0) <= NOT wire_y_pipeff_1_w_q_range865w(0);
	wire_y_pipeff_1_w_lg_w_q_range1033w1034w(0) <= NOT wire_y_pipeff_1_w_q_range1033w(0);
	wire_y_pipeff_1_w_lg_w_q_range1039w1040w(0) <= NOT wire_y_pipeff_1_w_q_range1039w(0);
	wire_y_pipeff_1_w_lg_w_q_range1045w1046w(0) <= NOT wire_y_pipeff_1_w_q_range1045w(0);
	wire_y_pipeff_1_w_lg_w_q_range845w846w(0) <= NOT wire_y_pipeff_1_w_q_range845w(0);
	wire_y_pipeff_1_w_lg_w_q_range871w872w(0) <= NOT wire_y_pipeff_1_w_q_range871w(0);
	wire_y_pipeff_1_w_lg_w_q_range877w878w(0) <= NOT wire_y_pipeff_1_w_q_range877w(0);
	wire_y_pipeff_1_w_lg_w_q_range883w884w(0) <= NOT wire_y_pipeff_1_w_q_range883w(0);
	wire_y_pipeff_1_w_lg_w_q_range889w890w(0) <= NOT wire_y_pipeff_1_w_q_range889w(0);
	wire_y_pipeff_1_w_lg_w_q_range895w896w(0) <= NOT wire_y_pipeff_1_w_q_range895w(0);
	wire_y_pipeff_1_w_lg_w_q_range901w902w(0) <= NOT wire_y_pipeff_1_w_q_range901w(0);
	wire_y_pipeff_1_w_lg_w_q_range907w908w(0) <= NOT wire_y_pipeff_1_w_q_range907w(0);
	wire_y_pipeff_1_w_q_range913w(0) <= y_pipeff_1(10);
	wire_y_pipeff_1_w_q_range919w(0) <= y_pipeff_1(11);
	wire_y_pipeff_1_w_q_range925w(0) <= y_pipeff_1(12);
	wire_y_pipeff_1_w_q_range931w(0) <= y_pipeff_1(13);
	wire_y_pipeff_1_w_q_range937w(0) <= y_pipeff_1(14);
	wire_y_pipeff_1_w_q_range943w(0) <= y_pipeff_1(15);
	wire_y_pipeff_1_w_q_range949w(0) <= y_pipeff_1(16);
	wire_y_pipeff_1_w_q_range955w(0) <= y_pipeff_1(17);
	wire_y_pipeff_1_w_q_range961w(0) <= y_pipeff_1(18);
	wire_y_pipeff_1_w_q_range967w(0) <= y_pipeff_1(19);
	wire_y_pipeff_1_w_q_range860w(0) <= y_pipeff_1(1);
	wire_y_pipeff_1_w_q_range973w(0) <= y_pipeff_1(20);
	wire_y_pipeff_1_w_q_range979w(0) <= y_pipeff_1(21);
	wire_y_pipeff_1_w_q_range985w(0) <= y_pipeff_1(22);
	wire_y_pipeff_1_w_q_range991w(0) <= y_pipeff_1(23);
	wire_y_pipeff_1_w_q_range997w(0) <= y_pipeff_1(24);
	wire_y_pipeff_1_w_q_range1003w(0) <= y_pipeff_1(25);
	wire_y_pipeff_1_w_q_range1009w(0) <= y_pipeff_1(26);
	wire_y_pipeff_1_w_q_range1015w(0) <= y_pipeff_1(27);
	wire_y_pipeff_1_w_q_range1021w(0) <= y_pipeff_1(28);
	wire_y_pipeff_1_w_q_range1027w(0) <= y_pipeff_1(29);
	wire_y_pipeff_1_w_q_range865w(0) <= y_pipeff_1(2);
	wire_y_pipeff_1_w_q_range1033w(0) <= y_pipeff_1(30);
	wire_y_pipeff_1_w_q_range1039w(0) <= y_pipeff_1(31);
	wire_y_pipeff_1_w_q_range1045w(0) <= y_pipeff_1(32);
	wire_y_pipeff_1_w_q_range845w(0) <= y_pipeff_1(33);
	wire_y_pipeff_1_w_q_range871w(0) <= y_pipeff_1(3);
	wire_y_pipeff_1_w_q_range877w(0) <= y_pipeff_1(4);
	wire_y_pipeff_1_w_q_range883w(0) <= y_pipeff_1(5);
	wire_y_pipeff_1_w_q_range889w(0) <= y_pipeff_1(6);
	wire_y_pipeff_1_w_q_range895w(0) <= y_pipeff_1(7);
	wire_y_pipeff_1_w_q_range901w(0) <= y_pipeff_1(8);
	wire_y_pipeff_1_w_q_range907w(0) <= y_pipeff_1(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_10 <= y_pipenode_10_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_10_w_lg_w_q_range8384w8385w(0) <= NOT wire_y_pipeff_10_w_q_range8384w(0);
	wire_y_pipeff_10_w_lg_w_q_range8389w8390w(0) <= NOT wire_y_pipeff_10_w_q_range8389w(0);
	wire_y_pipeff_10_w_lg_w_q_range8395w8396w(0) <= NOT wire_y_pipeff_10_w_q_range8395w(0);
	wire_y_pipeff_10_w_lg_w_q_range8401w8402w(0) <= NOT wire_y_pipeff_10_w_q_range8401w(0);
	wire_y_pipeff_10_w_lg_w_q_range8407w8408w(0) <= NOT wire_y_pipeff_10_w_q_range8407w(0);
	wire_y_pipeff_10_w_lg_w_q_range8413w8414w(0) <= NOT wire_y_pipeff_10_w_q_range8413w(0);
	wire_y_pipeff_10_w_lg_w_q_range8419w8420w(0) <= NOT wire_y_pipeff_10_w_q_range8419w(0);
	wire_y_pipeff_10_w_lg_w_q_range8425w8426w(0) <= NOT wire_y_pipeff_10_w_q_range8425w(0);
	wire_y_pipeff_10_w_lg_w_q_range8431w8432w(0) <= NOT wire_y_pipeff_10_w_q_range8431w(0);
	wire_y_pipeff_10_w_lg_w_q_range8437w8438w(0) <= NOT wire_y_pipeff_10_w_q_range8437w(0);
	wire_y_pipeff_10_w_lg_w_q_range8443w8444w(0) <= NOT wire_y_pipeff_10_w_q_range8443w(0);
	wire_y_pipeff_10_w_lg_w_q_range8449w8450w(0) <= NOT wire_y_pipeff_10_w_q_range8449w(0);
	wire_y_pipeff_10_w_lg_w_q_range8455w8456w(0) <= NOT wire_y_pipeff_10_w_q_range8455w(0);
	wire_y_pipeff_10_w_lg_w_q_range8461w8462w(0) <= NOT wire_y_pipeff_10_w_q_range8461w(0);
	wire_y_pipeff_10_w_lg_w_q_range8467w8468w(0) <= NOT wire_y_pipeff_10_w_q_range8467w(0);
	wire_y_pipeff_10_w_lg_w_q_range8473w8474w(0) <= NOT wire_y_pipeff_10_w_q_range8473w(0);
	wire_y_pipeff_10_w_lg_w_q_range8479w8480w(0) <= NOT wire_y_pipeff_10_w_q_range8479w(0);
	wire_y_pipeff_10_w_lg_w_q_range8485w8486w(0) <= NOT wire_y_pipeff_10_w_q_range8485w(0);
	wire_y_pipeff_10_w_lg_w_q_range8491w8492w(0) <= NOT wire_y_pipeff_10_w_q_range8491w(0);
	wire_y_pipeff_10_w_lg_w_q_range8497w8498w(0) <= NOT wire_y_pipeff_10_w_q_range8497w(0);
	wire_y_pipeff_10_w_lg_w_q_range8503w8504w(0) <= NOT wire_y_pipeff_10_w_q_range8503w(0);
	wire_y_pipeff_10_w_lg_w_q_range8509w8510w(0) <= NOT wire_y_pipeff_10_w_q_range8509w(0);
	wire_y_pipeff_10_w_lg_w_q_range8515w8516w(0) <= NOT wire_y_pipeff_10_w_q_range8515w(0);
	wire_y_pipeff_10_w_lg_w_q_range8333w8334w(0) <= NOT wire_y_pipeff_10_w_q_range8333w(0);
	wire_y_pipeff_10_w_q_range8384w(0) <= y_pipeff_10(10);
	wire_y_pipeff_10_w_q_range8389w(0) <= y_pipeff_10(11);
	wire_y_pipeff_10_w_q_range8395w(0) <= y_pipeff_10(12);
	wire_y_pipeff_10_w_q_range8401w(0) <= y_pipeff_10(13);
	wire_y_pipeff_10_w_q_range8407w(0) <= y_pipeff_10(14);
	wire_y_pipeff_10_w_q_range8413w(0) <= y_pipeff_10(15);
	wire_y_pipeff_10_w_q_range8419w(0) <= y_pipeff_10(16);
	wire_y_pipeff_10_w_q_range8425w(0) <= y_pipeff_10(17);
	wire_y_pipeff_10_w_q_range8431w(0) <= y_pipeff_10(18);
	wire_y_pipeff_10_w_q_range8437w(0) <= y_pipeff_10(19);
	wire_y_pipeff_10_w_q_range8443w(0) <= y_pipeff_10(20);
	wire_y_pipeff_10_w_q_range8449w(0) <= y_pipeff_10(21);
	wire_y_pipeff_10_w_q_range8455w(0) <= y_pipeff_10(22);
	wire_y_pipeff_10_w_q_range8461w(0) <= y_pipeff_10(23);
	wire_y_pipeff_10_w_q_range8467w(0) <= y_pipeff_10(24);
	wire_y_pipeff_10_w_q_range8473w(0) <= y_pipeff_10(25);
	wire_y_pipeff_10_w_q_range8479w(0) <= y_pipeff_10(26);
	wire_y_pipeff_10_w_q_range8485w(0) <= y_pipeff_10(27);
	wire_y_pipeff_10_w_q_range8491w(0) <= y_pipeff_10(28);
	wire_y_pipeff_10_w_q_range8497w(0) <= y_pipeff_10(29);
	wire_y_pipeff_10_w_q_range8503w(0) <= y_pipeff_10(30);
	wire_y_pipeff_10_w_q_range8509w(0) <= y_pipeff_10(31);
	wire_y_pipeff_10_w_q_range8515w(0) <= y_pipeff_10(32);
	wire_y_pipeff_10_w_q_range8333w(0) <= y_pipeff_10(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_11 <= y_pipenode_11_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_11_w_lg_w_q_range9195w9196w(0) <= NOT wire_y_pipeff_11_w_q_range9195w(0);
	wire_y_pipeff_11_w_lg_w_q_range9200w9201w(0) <= NOT wire_y_pipeff_11_w_q_range9200w(0);
	wire_y_pipeff_11_w_lg_w_q_range9206w9207w(0) <= NOT wire_y_pipeff_11_w_q_range9206w(0);
	wire_y_pipeff_11_w_lg_w_q_range9212w9213w(0) <= NOT wire_y_pipeff_11_w_q_range9212w(0);
	wire_y_pipeff_11_w_lg_w_q_range9218w9219w(0) <= NOT wire_y_pipeff_11_w_q_range9218w(0);
	wire_y_pipeff_11_w_lg_w_q_range9224w9225w(0) <= NOT wire_y_pipeff_11_w_q_range9224w(0);
	wire_y_pipeff_11_w_lg_w_q_range9230w9231w(0) <= NOT wire_y_pipeff_11_w_q_range9230w(0);
	wire_y_pipeff_11_w_lg_w_q_range9236w9237w(0) <= NOT wire_y_pipeff_11_w_q_range9236w(0);
	wire_y_pipeff_11_w_lg_w_q_range9242w9243w(0) <= NOT wire_y_pipeff_11_w_q_range9242w(0);
	wire_y_pipeff_11_w_lg_w_q_range9248w9249w(0) <= NOT wire_y_pipeff_11_w_q_range9248w(0);
	wire_y_pipeff_11_w_lg_w_q_range9254w9255w(0) <= NOT wire_y_pipeff_11_w_q_range9254w(0);
	wire_y_pipeff_11_w_lg_w_q_range9260w9261w(0) <= NOT wire_y_pipeff_11_w_q_range9260w(0);
	wire_y_pipeff_11_w_lg_w_q_range9266w9267w(0) <= NOT wire_y_pipeff_11_w_q_range9266w(0);
	wire_y_pipeff_11_w_lg_w_q_range9272w9273w(0) <= NOT wire_y_pipeff_11_w_q_range9272w(0);
	wire_y_pipeff_11_w_lg_w_q_range9278w9279w(0) <= NOT wire_y_pipeff_11_w_q_range9278w(0);
	wire_y_pipeff_11_w_lg_w_q_range9284w9285w(0) <= NOT wire_y_pipeff_11_w_q_range9284w(0);
	wire_y_pipeff_11_w_lg_w_q_range9290w9291w(0) <= NOT wire_y_pipeff_11_w_q_range9290w(0);
	wire_y_pipeff_11_w_lg_w_q_range9296w9297w(0) <= NOT wire_y_pipeff_11_w_q_range9296w(0);
	wire_y_pipeff_11_w_lg_w_q_range9302w9303w(0) <= NOT wire_y_pipeff_11_w_q_range9302w(0);
	wire_y_pipeff_11_w_lg_w_q_range9308w9309w(0) <= NOT wire_y_pipeff_11_w_q_range9308w(0);
	wire_y_pipeff_11_w_lg_w_q_range9314w9315w(0) <= NOT wire_y_pipeff_11_w_q_range9314w(0);
	wire_y_pipeff_11_w_lg_w_q_range9320w9321w(0) <= NOT wire_y_pipeff_11_w_q_range9320w(0);
	wire_y_pipeff_11_w_lg_w_q_range9140w9141w(0) <= NOT wire_y_pipeff_11_w_q_range9140w(0);
	wire_y_pipeff_11_w_q_range9195w(0) <= y_pipeff_11(11);
	wire_y_pipeff_11_w_q_range9200w(0) <= y_pipeff_11(12);
	wire_y_pipeff_11_w_q_range9206w(0) <= y_pipeff_11(13);
	wire_y_pipeff_11_w_q_range9212w(0) <= y_pipeff_11(14);
	wire_y_pipeff_11_w_q_range9218w(0) <= y_pipeff_11(15);
	wire_y_pipeff_11_w_q_range9224w(0) <= y_pipeff_11(16);
	wire_y_pipeff_11_w_q_range9230w(0) <= y_pipeff_11(17);
	wire_y_pipeff_11_w_q_range9236w(0) <= y_pipeff_11(18);
	wire_y_pipeff_11_w_q_range9242w(0) <= y_pipeff_11(19);
	wire_y_pipeff_11_w_q_range9248w(0) <= y_pipeff_11(20);
	wire_y_pipeff_11_w_q_range9254w(0) <= y_pipeff_11(21);
	wire_y_pipeff_11_w_q_range9260w(0) <= y_pipeff_11(22);
	wire_y_pipeff_11_w_q_range9266w(0) <= y_pipeff_11(23);
	wire_y_pipeff_11_w_q_range9272w(0) <= y_pipeff_11(24);
	wire_y_pipeff_11_w_q_range9278w(0) <= y_pipeff_11(25);
	wire_y_pipeff_11_w_q_range9284w(0) <= y_pipeff_11(26);
	wire_y_pipeff_11_w_q_range9290w(0) <= y_pipeff_11(27);
	wire_y_pipeff_11_w_q_range9296w(0) <= y_pipeff_11(28);
	wire_y_pipeff_11_w_q_range9302w(0) <= y_pipeff_11(29);
	wire_y_pipeff_11_w_q_range9308w(0) <= y_pipeff_11(30);
	wire_y_pipeff_11_w_q_range9314w(0) <= y_pipeff_11(31);
	wire_y_pipeff_11_w_q_range9320w(0) <= y_pipeff_11(32);
	wire_y_pipeff_11_w_q_range9140w(0) <= y_pipeff_11(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_12 <= y_pipenode_12_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_12_w_lg_w_q_range10001w10002w(0) <= NOT wire_y_pipeff_12_w_q_range10001w(0);
	wire_y_pipeff_12_w_lg_w_q_range10006w10007w(0) <= NOT wire_y_pipeff_12_w_q_range10006w(0);
	wire_y_pipeff_12_w_lg_w_q_range10012w10013w(0) <= NOT wire_y_pipeff_12_w_q_range10012w(0);
	wire_y_pipeff_12_w_lg_w_q_range10018w10019w(0) <= NOT wire_y_pipeff_12_w_q_range10018w(0);
	wire_y_pipeff_12_w_lg_w_q_range10024w10025w(0) <= NOT wire_y_pipeff_12_w_q_range10024w(0);
	wire_y_pipeff_12_w_lg_w_q_range10030w10031w(0) <= NOT wire_y_pipeff_12_w_q_range10030w(0);
	wire_y_pipeff_12_w_lg_w_q_range10036w10037w(0) <= NOT wire_y_pipeff_12_w_q_range10036w(0);
	wire_y_pipeff_12_w_lg_w_q_range10042w10043w(0) <= NOT wire_y_pipeff_12_w_q_range10042w(0);
	wire_y_pipeff_12_w_lg_w_q_range10048w10049w(0) <= NOT wire_y_pipeff_12_w_q_range10048w(0);
	wire_y_pipeff_12_w_lg_w_q_range10054w10055w(0) <= NOT wire_y_pipeff_12_w_q_range10054w(0);
	wire_y_pipeff_12_w_lg_w_q_range10060w10061w(0) <= NOT wire_y_pipeff_12_w_q_range10060w(0);
	wire_y_pipeff_12_w_lg_w_q_range10066w10067w(0) <= NOT wire_y_pipeff_12_w_q_range10066w(0);
	wire_y_pipeff_12_w_lg_w_q_range10072w10073w(0) <= NOT wire_y_pipeff_12_w_q_range10072w(0);
	wire_y_pipeff_12_w_lg_w_q_range10078w10079w(0) <= NOT wire_y_pipeff_12_w_q_range10078w(0);
	wire_y_pipeff_12_w_lg_w_q_range10084w10085w(0) <= NOT wire_y_pipeff_12_w_q_range10084w(0);
	wire_y_pipeff_12_w_lg_w_q_range10090w10091w(0) <= NOT wire_y_pipeff_12_w_q_range10090w(0);
	wire_y_pipeff_12_w_lg_w_q_range10096w10097w(0) <= NOT wire_y_pipeff_12_w_q_range10096w(0);
	wire_y_pipeff_12_w_lg_w_q_range10102w10103w(0) <= NOT wire_y_pipeff_12_w_q_range10102w(0);
	wire_y_pipeff_12_w_lg_w_q_range10108w10109w(0) <= NOT wire_y_pipeff_12_w_q_range10108w(0);
	wire_y_pipeff_12_w_lg_w_q_range10114w10115w(0) <= NOT wire_y_pipeff_12_w_q_range10114w(0);
	wire_y_pipeff_12_w_lg_w_q_range10120w10121w(0) <= NOT wire_y_pipeff_12_w_q_range10120w(0);
	wire_y_pipeff_12_w_lg_w_q_range9942w9943w(0) <= NOT wire_y_pipeff_12_w_q_range9942w(0);
	wire_y_pipeff_12_w_q_range10001w(0) <= y_pipeff_12(12);
	wire_y_pipeff_12_w_q_range10006w(0) <= y_pipeff_12(13);
	wire_y_pipeff_12_w_q_range10012w(0) <= y_pipeff_12(14);
	wire_y_pipeff_12_w_q_range10018w(0) <= y_pipeff_12(15);
	wire_y_pipeff_12_w_q_range10024w(0) <= y_pipeff_12(16);
	wire_y_pipeff_12_w_q_range10030w(0) <= y_pipeff_12(17);
	wire_y_pipeff_12_w_q_range10036w(0) <= y_pipeff_12(18);
	wire_y_pipeff_12_w_q_range10042w(0) <= y_pipeff_12(19);
	wire_y_pipeff_12_w_q_range10048w(0) <= y_pipeff_12(20);
	wire_y_pipeff_12_w_q_range10054w(0) <= y_pipeff_12(21);
	wire_y_pipeff_12_w_q_range10060w(0) <= y_pipeff_12(22);
	wire_y_pipeff_12_w_q_range10066w(0) <= y_pipeff_12(23);
	wire_y_pipeff_12_w_q_range10072w(0) <= y_pipeff_12(24);
	wire_y_pipeff_12_w_q_range10078w(0) <= y_pipeff_12(25);
	wire_y_pipeff_12_w_q_range10084w(0) <= y_pipeff_12(26);
	wire_y_pipeff_12_w_q_range10090w(0) <= y_pipeff_12(27);
	wire_y_pipeff_12_w_q_range10096w(0) <= y_pipeff_12(28);
	wire_y_pipeff_12_w_q_range10102w(0) <= y_pipeff_12(29);
	wire_y_pipeff_12_w_q_range10108w(0) <= y_pipeff_12(30);
	wire_y_pipeff_12_w_q_range10114w(0) <= y_pipeff_12(31);
	wire_y_pipeff_12_w_q_range10120w(0) <= y_pipeff_12(32);
	wire_y_pipeff_12_w_q_range9942w(0) <= y_pipeff_12(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_13 <= y_pipenode_13_w;
			END IF;
		END IF;
	END PROCESS;
	loop34 : FOR i IN 0 TO 33 GENERATE 
		wire_y_pipeff_13_w_lg_q10740w(i) <= y_pipeff_13(i) AND wire_sincosbitff_w_lg_w_q_range668w10739w(0);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 33 GENERATE 
		wire_y_pipeff_13_w_lg_q10743w(i) <= y_pipeff_13(i) AND wire_sincosbitff_w_q_range668w(0);
	END GENERATE loop35;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_2 <= y_pipenode_2_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_2_w_lg_w_q_range1763w1764w(0) <= NOT wire_y_pipeff_2_w_q_range1763w(0);
	wire_y_pipeff_2_w_lg_w_q_range1769w1770w(0) <= NOT wire_y_pipeff_2_w_q_range1769w(0);
	wire_y_pipeff_2_w_lg_w_q_range1775w1776w(0) <= NOT wire_y_pipeff_2_w_q_range1775w(0);
	wire_y_pipeff_2_w_lg_w_q_range1781w1782w(0) <= NOT wire_y_pipeff_2_w_q_range1781w(0);
	wire_y_pipeff_2_w_lg_w_q_range1787w1788w(0) <= NOT wire_y_pipeff_2_w_q_range1787w(0);
	wire_y_pipeff_2_w_lg_w_q_range1793w1794w(0) <= NOT wire_y_pipeff_2_w_q_range1793w(0);
	wire_y_pipeff_2_w_lg_w_q_range1799w1800w(0) <= NOT wire_y_pipeff_2_w_q_range1799w(0);
	wire_y_pipeff_2_w_lg_w_q_range1805w1806w(0) <= NOT wire_y_pipeff_2_w_q_range1805w(0);
	wire_y_pipeff_2_w_lg_w_q_range1811w1812w(0) <= NOT wire_y_pipeff_2_w_q_range1811w(0);
	wire_y_pipeff_2_w_lg_w_q_range1817w1818w(0) <= NOT wire_y_pipeff_2_w_q_range1817w(0);
	wire_y_pipeff_2_w_lg_w_q_range1823w1824w(0) <= NOT wire_y_pipeff_2_w_q_range1823w(0);
	wire_y_pipeff_2_w_lg_w_q_range1829w1830w(0) <= NOT wire_y_pipeff_2_w_q_range1829w(0);
	wire_y_pipeff_2_w_lg_w_q_range1835w1836w(0) <= NOT wire_y_pipeff_2_w_q_range1835w(0);
	wire_y_pipeff_2_w_lg_w_q_range1841w1842w(0) <= NOT wire_y_pipeff_2_w_q_range1841w(0);
	wire_y_pipeff_2_w_lg_w_q_range1847w1848w(0) <= NOT wire_y_pipeff_2_w_q_range1847w(0);
	wire_y_pipeff_2_w_lg_w_q_range1853w1854w(0) <= NOT wire_y_pipeff_2_w_q_range1853w(0);
	wire_y_pipeff_2_w_lg_w_q_range1859w1860w(0) <= NOT wire_y_pipeff_2_w_q_range1859w(0);
	wire_y_pipeff_2_w_lg_w_q_range1865w1866w(0) <= NOT wire_y_pipeff_2_w_q_range1865w(0);
	wire_y_pipeff_2_w_lg_w_q_range1871w1872w(0) <= NOT wire_y_pipeff_2_w_q_range1871w(0);
	wire_y_pipeff_2_w_lg_w_q_range1877w1878w(0) <= NOT wire_y_pipeff_2_w_q_range1877w(0);
	wire_y_pipeff_2_w_lg_w_q_range1716w1717w(0) <= NOT wire_y_pipeff_2_w_q_range1716w(0);
	wire_y_pipeff_2_w_lg_w_q_range1883w1884w(0) <= NOT wire_y_pipeff_2_w_q_range1883w(0);
	wire_y_pipeff_2_w_lg_w_q_range1889w1890w(0) <= NOT wire_y_pipeff_2_w_q_range1889w(0);
	wire_y_pipeff_2_w_lg_w_q_range1895w1896w(0) <= NOT wire_y_pipeff_2_w_q_range1895w(0);
	wire_y_pipeff_2_w_lg_w_q_range1697w1698w(0) <= NOT wire_y_pipeff_2_w_q_range1697w(0);
	wire_y_pipeff_2_w_lg_w_q_range1721w1722w(0) <= NOT wire_y_pipeff_2_w_q_range1721w(0);
	wire_y_pipeff_2_w_lg_w_q_range1727w1728w(0) <= NOT wire_y_pipeff_2_w_q_range1727w(0);
	wire_y_pipeff_2_w_lg_w_q_range1733w1734w(0) <= NOT wire_y_pipeff_2_w_q_range1733w(0);
	wire_y_pipeff_2_w_lg_w_q_range1739w1740w(0) <= NOT wire_y_pipeff_2_w_q_range1739w(0);
	wire_y_pipeff_2_w_lg_w_q_range1745w1746w(0) <= NOT wire_y_pipeff_2_w_q_range1745w(0);
	wire_y_pipeff_2_w_lg_w_q_range1751w1752w(0) <= NOT wire_y_pipeff_2_w_q_range1751w(0);
	wire_y_pipeff_2_w_lg_w_q_range1757w1758w(0) <= NOT wire_y_pipeff_2_w_q_range1757w(0);
	wire_y_pipeff_2_w_q_range1763w(0) <= y_pipeff_2(10);
	wire_y_pipeff_2_w_q_range1769w(0) <= y_pipeff_2(11);
	wire_y_pipeff_2_w_q_range1775w(0) <= y_pipeff_2(12);
	wire_y_pipeff_2_w_q_range1781w(0) <= y_pipeff_2(13);
	wire_y_pipeff_2_w_q_range1787w(0) <= y_pipeff_2(14);
	wire_y_pipeff_2_w_q_range1793w(0) <= y_pipeff_2(15);
	wire_y_pipeff_2_w_q_range1799w(0) <= y_pipeff_2(16);
	wire_y_pipeff_2_w_q_range1805w(0) <= y_pipeff_2(17);
	wire_y_pipeff_2_w_q_range1811w(0) <= y_pipeff_2(18);
	wire_y_pipeff_2_w_q_range1817w(0) <= y_pipeff_2(19);
	wire_y_pipeff_2_w_q_range1823w(0) <= y_pipeff_2(20);
	wire_y_pipeff_2_w_q_range1829w(0) <= y_pipeff_2(21);
	wire_y_pipeff_2_w_q_range1835w(0) <= y_pipeff_2(22);
	wire_y_pipeff_2_w_q_range1841w(0) <= y_pipeff_2(23);
	wire_y_pipeff_2_w_q_range1847w(0) <= y_pipeff_2(24);
	wire_y_pipeff_2_w_q_range1853w(0) <= y_pipeff_2(25);
	wire_y_pipeff_2_w_q_range1859w(0) <= y_pipeff_2(26);
	wire_y_pipeff_2_w_q_range1865w(0) <= y_pipeff_2(27);
	wire_y_pipeff_2_w_q_range1871w(0) <= y_pipeff_2(28);
	wire_y_pipeff_2_w_q_range1877w(0) <= y_pipeff_2(29);
	wire_y_pipeff_2_w_q_range1716w(0) <= y_pipeff_2(2);
	wire_y_pipeff_2_w_q_range1883w(0) <= y_pipeff_2(30);
	wire_y_pipeff_2_w_q_range1889w(0) <= y_pipeff_2(31);
	wire_y_pipeff_2_w_q_range1895w(0) <= y_pipeff_2(32);
	wire_y_pipeff_2_w_q_range1697w(0) <= y_pipeff_2(33);
	wire_y_pipeff_2_w_q_range1721w(0) <= y_pipeff_2(3);
	wire_y_pipeff_2_w_q_range1727w(0) <= y_pipeff_2(4);
	wire_y_pipeff_2_w_q_range1733w(0) <= y_pipeff_2(5);
	wire_y_pipeff_2_w_q_range1739w(0) <= y_pipeff_2(6);
	wire_y_pipeff_2_w_q_range1745w(0) <= y_pipeff_2(7);
	wire_y_pipeff_2_w_q_range1751w(0) <= y_pipeff_2(8);
	wire_y_pipeff_2_w_q_range1757w(0) <= y_pipeff_2(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_3 <= y_pipenode_3_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_3_w_lg_w_q_range2608w2609w(0) <= NOT wire_y_pipeff_3_w_q_range2608w(0);
	wire_y_pipeff_3_w_lg_w_q_range2614w2615w(0) <= NOT wire_y_pipeff_3_w_q_range2614w(0);
	wire_y_pipeff_3_w_lg_w_q_range2620w2621w(0) <= NOT wire_y_pipeff_3_w_q_range2620w(0);
	wire_y_pipeff_3_w_lg_w_q_range2626w2627w(0) <= NOT wire_y_pipeff_3_w_q_range2626w(0);
	wire_y_pipeff_3_w_lg_w_q_range2632w2633w(0) <= NOT wire_y_pipeff_3_w_q_range2632w(0);
	wire_y_pipeff_3_w_lg_w_q_range2638w2639w(0) <= NOT wire_y_pipeff_3_w_q_range2638w(0);
	wire_y_pipeff_3_w_lg_w_q_range2644w2645w(0) <= NOT wire_y_pipeff_3_w_q_range2644w(0);
	wire_y_pipeff_3_w_lg_w_q_range2650w2651w(0) <= NOT wire_y_pipeff_3_w_q_range2650w(0);
	wire_y_pipeff_3_w_lg_w_q_range2656w2657w(0) <= NOT wire_y_pipeff_3_w_q_range2656w(0);
	wire_y_pipeff_3_w_lg_w_q_range2662w2663w(0) <= NOT wire_y_pipeff_3_w_q_range2662w(0);
	wire_y_pipeff_3_w_lg_w_q_range2668w2669w(0) <= NOT wire_y_pipeff_3_w_q_range2668w(0);
	wire_y_pipeff_3_w_lg_w_q_range2674w2675w(0) <= NOT wire_y_pipeff_3_w_q_range2674w(0);
	wire_y_pipeff_3_w_lg_w_q_range2680w2681w(0) <= NOT wire_y_pipeff_3_w_q_range2680w(0);
	wire_y_pipeff_3_w_lg_w_q_range2686w2687w(0) <= NOT wire_y_pipeff_3_w_q_range2686w(0);
	wire_y_pipeff_3_w_lg_w_q_range2692w2693w(0) <= NOT wire_y_pipeff_3_w_q_range2692w(0);
	wire_y_pipeff_3_w_lg_w_q_range2698w2699w(0) <= NOT wire_y_pipeff_3_w_q_range2698w(0);
	wire_y_pipeff_3_w_lg_w_q_range2704w2705w(0) <= NOT wire_y_pipeff_3_w_q_range2704w(0);
	wire_y_pipeff_3_w_lg_w_q_range2710w2711w(0) <= NOT wire_y_pipeff_3_w_q_range2710w(0);
	wire_y_pipeff_3_w_lg_w_q_range2716w2717w(0) <= NOT wire_y_pipeff_3_w_q_range2716w(0);
	wire_y_pipeff_3_w_lg_w_q_range2722w2723w(0) <= NOT wire_y_pipeff_3_w_q_range2722w(0);
	wire_y_pipeff_3_w_lg_w_q_range2728w2729w(0) <= NOT wire_y_pipeff_3_w_q_range2728w(0);
	wire_y_pipeff_3_w_lg_w_q_range2734w2735w(0) <= NOT wire_y_pipeff_3_w_q_range2734w(0);
	wire_y_pipeff_3_w_lg_w_q_range2740w2741w(0) <= NOT wire_y_pipeff_3_w_q_range2740w(0);
	wire_y_pipeff_3_w_lg_w_q_range2544w2545w(0) <= NOT wire_y_pipeff_3_w_q_range2544w(0);
	wire_y_pipeff_3_w_lg_w_q_range2567w2568w(0) <= NOT wire_y_pipeff_3_w_q_range2567w(0);
	wire_y_pipeff_3_w_lg_w_q_range2572w2573w(0) <= NOT wire_y_pipeff_3_w_q_range2572w(0);
	wire_y_pipeff_3_w_lg_w_q_range2578w2579w(0) <= NOT wire_y_pipeff_3_w_q_range2578w(0);
	wire_y_pipeff_3_w_lg_w_q_range2584w2585w(0) <= NOT wire_y_pipeff_3_w_q_range2584w(0);
	wire_y_pipeff_3_w_lg_w_q_range2590w2591w(0) <= NOT wire_y_pipeff_3_w_q_range2590w(0);
	wire_y_pipeff_3_w_lg_w_q_range2596w2597w(0) <= NOT wire_y_pipeff_3_w_q_range2596w(0);
	wire_y_pipeff_3_w_lg_w_q_range2602w2603w(0) <= NOT wire_y_pipeff_3_w_q_range2602w(0);
	wire_y_pipeff_3_w_q_range2608w(0) <= y_pipeff_3(10);
	wire_y_pipeff_3_w_q_range2614w(0) <= y_pipeff_3(11);
	wire_y_pipeff_3_w_q_range2620w(0) <= y_pipeff_3(12);
	wire_y_pipeff_3_w_q_range2626w(0) <= y_pipeff_3(13);
	wire_y_pipeff_3_w_q_range2632w(0) <= y_pipeff_3(14);
	wire_y_pipeff_3_w_q_range2638w(0) <= y_pipeff_3(15);
	wire_y_pipeff_3_w_q_range2644w(0) <= y_pipeff_3(16);
	wire_y_pipeff_3_w_q_range2650w(0) <= y_pipeff_3(17);
	wire_y_pipeff_3_w_q_range2656w(0) <= y_pipeff_3(18);
	wire_y_pipeff_3_w_q_range2662w(0) <= y_pipeff_3(19);
	wire_y_pipeff_3_w_q_range2668w(0) <= y_pipeff_3(20);
	wire_y_pipeff_3_w_q_range2674w(0) <= y_pipeff_3(21);
	wire_y_pipeff_3_w_q_range2680w(0) <= y_pipeff_3(22);
	wire_y_pipeff_3_w_q_range2686w(0) <= y_pipeff_3(23);
	wire_y_pipeff_3_w_q_range2692w(0) <= y_pipeff_3(24);
	wire_y_pipeff_3_w_q_range2698w(0) <= y_pipeff_3(25);
	wire_y_pipeff_3_w_q_range2704w(0) <= y_pipeff_3(26);
	wire_y_pipeff_3_w_q_range2710w(0) <= y_pipeff_3(27);
	wire_y_pipeff_3_w_q_range2716w(0) <= y_pipeff_3(28);
	wire_y_pipeff_3_w_q_range2722w(0) <= y_pipeff_3(29);
	wire_y_pipeff_3_w_q_range2728w(0) <= y_pipeff_3(30);
	wire_y_pipeff_3_w_q_range2734w(0) <= y_pipeff_3(31);
	wire_y_pipeff_3_w_q_range2740w(0) <= y_pipeff_3(32);
	wire_y_pipeff_3_w_q_range2544w(0) <= y_pipeff_3(33);
	wire_y_pipeff_3_w_q_range2567w(0) <= y_pipeff_3(3);
	wire_y_pipeff_3_w_q_range2572w(0) <= y_pipeff_3(4);
	wire_y_pipeff_3_w_q_range2578w(0) <= y_pipeff_3(5);
	wire_y_pipeff_3_w_q_range2584w(0) <= y_pipeff_3(6);
	wire_y_pipeff_3_w_q_range2590w(0) <= y_pipeff_3(7);
	wire_y_pipeff_3_w_q_range2596w(0) <= y_pipeff_3(8);
	wire_y_pipeff_3_w_q_range2602w(0) <= y_pipeff_3(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_4 <= y_pipenode_4_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_4_w_lg_w_q_range3448w3449w(0) <= NOT wire_y_pipeff_4_w_q_range3448w(0);
	wire_y_pipeff_4_w_lg_w_q_range3454w3455w(0) <= NOT wire_y_pipeff_4_w_q_range3454w(0);
	wire_y_pipeff_4_w_lg_w_q_range3460w3461w(0) <= NOT wire_y_pipeff_4_w_q_range3460w(0);
	wire_y_pipeff_4_w_lg_w_q_range3466w3467w(0) <= NOT wire_y_pipeff_4_w_q_range3466w(0);
	wire_y_pipeff_4_w_lg_w_q_range3472w3473w(0) <= NOT wire_y_pipeff_4_w_q_range3472w(0);
	wire_y_pipeff_4_w_lg_w_q_range3478w3479w(0) <= NOT wire_y_pipeff_4_w_q_range3478w(0);
	wire_y_pipeff_4_w_lg_w_q_range3484w3485w(0) <= NOT wire_y_pipeff_4_w_q_range3484w(0);
	wire_y_pipeff_4_w_lg_w_q_range3490w3491w(0) <= NOT wire_y_pipeff_4_w_q_range3490w(0);
	wire_y_pipeff_4_w_lg_w_q_range3496w3497w(0) <= NOT wire_y_pipeff_4_w_q_range3496w(0);
	wire_y_pipeff_4_w_lg_w_q_range3502w3503w(0) <= NOT wire_y_pipeff_4_w_q_range3502w(0);
	wire_y_pipeff_4_w_lg_w_q_range3508w3509w(0) <= NOT wire_y_pipeff_4_w_q_range3508w(0);
	wire_y_pipeff_4_w_lg_w_q_range3514w3515w(0) <= NOT wire_y_pipeff_4_w_q_range3514w(0);
	wire_y_pipeff_4_w_lg_w_q_range3520w3521w(0) <= NOT wire_y_pipeff_4_w_q_range3520w(0);
	wire_y_pipeff_4_w_lg_w_q_range3526w3527w(0) <= NOT wire_y_pipeff_4_w_q_range3526w(0);
	wire_y_pipeff_4_w_lg_w_q_range3532w3533w(0) <= NOT wire_y_pipeff_4_w_q_range3532w(0);
	wire_y_pipeff_4_w_lg_w_q_range3538w3539w(0) <= NOT wire_y_pipeff_4_w_q_range3538w(0);
	wire_y_pipeff_4_w_lg_w_q_range3544w3545w(0) <= NOT wire_y_pipeff_4_w_q_range3544w(0);
	wire_y_pipeff_4_w_lg_w_q_range3550w3551w(0) <= NOT wire_y_pipeff_4_w_q_range3550w(0);
	wire_y_pipeff_4_w_lg_w_q_range3556w3557w(0) <= NOT wire_y_pipeff_4_w_q_range3556w(0);
	wire_y_pipeff_4_w_lg_w_q_range3562w3563w(0) <= NOT wire_y_pipeff_4_w_q_range3562w(0);
	wire_y_pipeff_4_w_lg_w_q_range3568w3569w(0) <= NOT wire_y_pipeff_4_w_q_range3568w(0);
	wire_y_pipeff_4_w_lg_w_q_range3574w3575w(0) <= NOT wire_y_pipeff_4_w_q_range3574w(0);
	wire_y_pipeff_4_w_lg_w_q_range3580w3581w(0) <= NOT wire_y_pipeff_4_w_q_range3580w(0);
	wire_y_pipeff_4_w_lg_w_q_range3386w3387w(0) <= NOT wire_y_pipeff_4_w_q_range3386w(0);
	wire_y_pipeff_4_w_lg_w_q_range3413w3414w(0) <= NOT wire_y_pipeff_4_w_q_range3413w(0);
	wire_y_pipeff_4_w_lg_w_q_range3418w3419w(0) <= NOT wire_y_pipeff_4_w_q_range3418w(0);
	wire_y_pipeff_4_w_lg_w_q_range3424w3425w(0) <= NOT wire_y_pipeff_4_w_q_range3424w(0);
	wire_y_pipeff_4_w_lg_w_q_range3430w3431w(0) <= NOT wire_y_pipeff_4_w_q_range3430w(0);
	wire_y_pipeff_4_w_lg_w_q_range3436w3437w(0) <= NOT wire_y_pipeff_4_w_q_range3436w(0);
	wire_y_pipeff_4_w_lg_w_q_range3442w3443w(0) <= NOT wire_y_pipeff_4_w_q_range3442w(0);
	wire_y_pipeff_4_w_q_range3448w(0) <= y_pipeff_4(10);
	wire_y_pipeff_4_w_q_range3454w(0) <= y_pipeff_4(11);
	wire_y_pipeff_4_w_q_range3460w(0) <= y_pipeff_4(12);
	wire_y_pipeff_4_w_q_range3466w(0) <= y_pipeff_4(13);
	wire_y_pipeff_4_w_q_range3472w(0) <= y_pipeff_4(14);
	wire_y_pipeff_4_w_q_range3478w(0) <= y_pipeff_4(15);
	wire_y_pipeff_4_w_q_range3484w(0) <= y_pipeff_4(16);
	wire_y_pipeff_4_w_q_range3490w(0) <= y_pipeff_4(17);
	wire_y_pipeff_4_w_q_range3496w(0) <= y_pipeff_4(18);
	wire_y_pipeff_4_w_q_range3502w(0) <= y_pipeff_4(19);
	wire_y_pipeff_4_w_q_range3508w(0) <= y_pipeff_4(20);
	wire_y_pipeff_4_w_q_range3514w(0) <= y_pipeff_4(21);
	wire_y_pipeff_4_w_q_range3520w(0) <= y_pipeff_4(22);
	wire_y_pipeff_4_w_q_range3526w(0) <= y_pipeff_4(23);
	wire_y_pipeff_4_w_q_range3532w(0) <= y_pipeff_4(24);
	wire_y_pipeff_4_w_q_range3538w(0) <= y_pipeff_4(25);
	wire_y_pipeff_4_w_q_range3544w(0) <= y_pipeff_4(26);
	wire_y_pipeff_4_w_q_range3550w(0) <= y_pipeff_4(27);
	wire_y_pipeff_4_w_q_range3556w(0) <= y_pipeff_4(28);
	wire_y_pipeff_4_w_q_range3562w(0) <= y_pipeff_4(29);
	wire_y_pipeff_4_w_q_range3568w(0) <= y_pipeff_4(30);
	wire_y_pipeff_4_w_q_range3574w(0) <= y_pipeff_4(31);
	wire_y_pipeff_4_w_q_range3580w(0) <= y_pipeff_4(32);
	wire_y_pipeff_4_w_q_range3386w(0) <= y_pipeff_4(33);
	wire_y_pipeff_4_w_q_range3413w(0) <= y_pipeff_4(4);
	wire_y_pipeff_4_w_q_range3418w(0) <= y_pipeff_4(5);
	wire_y_pipeff_4_w_q_range3424w(0) <= y_pipeff_4(6);
	wire_y_pipeff_4_w_q_range3430w(0) <= y_pipeff_4(7);
	wire_y_pipeff_4_w_q_range3436w(0) <= y_pipeff_4(8);
	wire_y_pipeff_4_w_q_range3442w(0) <= y_pipeff_4(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_5 <= y_pipenode_5_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_5_w_lg_w_q_range4283w4284w(0) <= NOT wire_y_pipeff_5_w_q_range4283w(0);
	wire_y_pipeff_5_w_lg_w_q_range4289w4290w(0) <= NOT wire_y_pipeff_5_w_q_range4289w(0);
	wire_y_pipeff_5_w_lg_w_q_range4295w4296w(0) <= NOT wire_y_pipeff_5_w_q_range4295w(0);
	wire_y_pipeff_5_w_lg_w_q_range4301w4302w(0) <= NOT wire_y_pipeff_5_w_q_range4301w(0);
	wire_y_pipeff_5_w_lg_w_q_range4307w4308w(0) <= NOT wire_y_pipeff_5_w_q_range4307w(0);
	wire_y_pipeff_5_w_lg_w_q_range4313w4314w(0) <= NOT wire_y_pipeff_5_w_q_range4313w(0);
	wire_y_pipeff_5_w_lg_w_q_range4319w4320w(0) <= NOT wire_y_pipeff_5_w_q_range4319w(0);
	wire_y_pipeff_5_w_lg_w_q_range4325w4326w(0) <= NOT wire_y_pipeff_5_w_q_range4325w(0);
	wire_y_pipeff_5_w_lg_w_q_range4331w4332w(0) <= NOT wire_y_pipeff_5_w_q_range4331w(0);
	wire_y_pipeff_5_w_lg_w_q_range4337w4338w(0) <= NOT wire_y_pipeff_5_w_q_range4337w(0);
	wire_y_pipeff_5_w_lg_w_q_range4343w4344w(0) <= NOT wire_y_pipeff_5_w_q_range4343w(0);
	wire_y_pipeff_5_w_lg_w_q_range4349w4350w(0) <= NOT wire_y_pipeff_5_w_q_range4349w(0);
	wire_y_pipeff_5_w_lg_w_q_range4355w4356w(0) <= NOT wire_y_pipeff_5_w_q_range4355w(0);
	wire_y_pipeff_5_w_lg_w_q_range4361w4362w(0) <= NOT wire_y_pipeff_5_w_q_range4361w(0);
	wire_y_pipeff_5_w_lg_w_q_range4367w4368w(0) <= NOT wire_y_pipeff_5_w_q_range4367w(0);
	wire_y_pipeff_5_w_lg_w_q_range4373w4374w(0) <= NOT wire_y_pipeff_5_w_q_range4373w(0);
	wire_y_pipeff_5_w_lg_w_q_range4379w4380w(0) <= NOT wire_y_pipeff_5_w_q_range4379w(0);
	wire_y_pipeff_5_w_lg_w_q_range4385w4386w(0) <= NOT wire_y_pipeff_5_w_q_range4385w(0);
	wire_y_pipeff_5_w_lg_w_q_range4391w4392w(0) <= NOT wire_y_pipeff_5_w_q_range4391w(0);
	wire_y_pipeff_5_w_lg_w_q_range4397w4398w(0) <= NOT wire_y_pipeff_5_w_q_range4397w(0);
	wire_y_pipeff_5_w_lg_w_q_range4403w4404w(0) <= NOT wire_y_pipeff_5_w_q_range4403w(0);
	wire_y_pipeff_5_w_lg_w_q_range4409w4410w(0) <= NOT wire_y_pipeff_5_w_q_range4409w(0);
	wire_y_pipeff_5_w_lg_w_q_range4415w4416w(0) <= NOT wire_y_pipeff_5_w_q_range4415w(0);
	wire_y_pipeff_5_w_lg_w_q_range4223w4224w(0) <= NOT wire_y_pipeff_5_w_q_range4223w(0);
	wire_y_pipeff_5_w_lg_w_q_range4254w4255w(0) <= NOT wire_y_pipeff_5_w_q_range4254w(0);
	wire_y_pipeff_5_w_lg_w_q_range4259w4260w(0) <= NOT wire_y_pipeff_5_w_q_range4259w(0);
	wire_y_pipeff_5_w_lg_w_q_range4265w4266w(0) <= NOT wire_y_pipeff_5_w_q_range4265w(0);
	wire_y_pipeff_5_w_lg_w_q_range4271w4272w(0) <= NOT wire_y_pipeff_5_w_q_range4271w(0);
	wire_y_pipeff_5_w_lg_w_q_range4277w4278w(0) <= NOT wire_y_pipeff_5_w_q_range4277w(0);
	wire_y_pipeff_5_w_q_range4283w(0) <= y_pipeff_5(10);
	wire_y_pipeff_5_w_q_range4289w(0) <= y_pipeff_5(11);
	wire_y_pipeff_5_w_q_range4295w(0) <= y_pipeff_5(12);
	wire_y_pipeff_5_w_q_range4301w(0) <= y_pipeff_5(13);
	wire_y_pipeff_5_w_q_range4307w(0) <= y_pipeff_5(14);
	wire_y_pipeff_5_w_q_range4313w(0) <= y_pipeff_5(15);
	wire_y_pipeff_5_w_q_range4319w(0) <= y_pipeff_5(16);
	wire_y_pipeff_5_w_q_range4325w(0) <= y_pipeff_5(17);
	wire_y_pipeff_5_w_q_range4331w(0) <= y_pipeff_5(18);
	wire_y_pipeff_5_w_q_range4337w(0) <= y_pipeff_5(19);
	wire_y_pipeff_5_w_q_range4343w(0) <= y_pipeff_5(20);
	wire_y_pipeff_5_w_q_range4349w(0) <= y_pipeff_5(21);
	wire_y_pipeff_5_w_q_range4355w(0) <= y_pipeff_5(22);
	wire_y_pipeff_5_w_q_range4361w(0) <= y_pipeff_5(23);
	wire_y_pipeff_5_w_q_range4367w(0) <= y_pipeff_5(24);
	wire_y_pipeff_5_w_q_range4373w(0) <= y_pipeff_5(25);
	wire_y_pipeff_5_w_q_range4379w(0) <= y_pipeff_5(26);
	wire_y_pipeff_5_w_q_range4385w(0) <= y_pipeff_5(27);
	wire_y_pipeff_5_w_q_range4391w(0) <= y_pipeff_5(28);
	wire_y_pipeff_5_w_q_range4397w(0) <= y_pipeff_5(29);
	wire_y_pipeff_5_w_q_range4403w(0) <= y_pipeff_5(30);
	wire_y_pipeff_5_w_q_range4409w(0) <= y_pipeff_5(31);
	wire_y_pipeff_5_w_q_range4415w(0) <= y_pipeff_5(32);
	wire_y_pipeff_5_w_q_range4223w(0) <= y_pipeff_5(33);
	wire_y_pipeff_5_w_q_range4254w(0) <= y_pipeff_5(5);
	wire_y_pipeff_5_w_q_range4259w(0) <= y_pipeff_5(6);
	wire_y_pipeff_5_w_q_range4265w(0) <= y_pipeff_5(7);
	wire_y_pipeff_5_w_q_range4271w(0) <= y_pipeff_5(8);
	wire_y_pipeff_5_w_q_range4277w(0) <= y_pipeff_5(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_6 <= y_pipenode_6_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_6_w_lg_w_q_range5113w5114w(0) <= NOT wire_y_pipeff_6_w_q_range5113w(0);
	wire_y_pipeff_6_w_lg_w_q_range5119w5120w(0) <= NOT wire_y_pipeff_6_w_q_range5119w(0);
	wire_y_pipeff_6_w_lg_w_q_range5125w5126w(0) <= NOT wire_y_pipeff_6_w_q_range5125w(0);
	wire_y_pipeff_6_w_lg_w_q_range5131w5132w(0) <= NOT wire_y_pipeff_6_w_q_range5131w(0);
	wire_y_pipeff_6_w_lg_w_q_range5137w5138w(0) <= NOT wire_y_pipeff_6_w_q_range5137w(0);
	wire_y_pipeff_6_w_lg_w_q_range5143w5144w(0) <= NOT wire_y_pipeff_6_w_q_range5143w(0);
	wire_y_pipeff_6_w_lg_w_q_range5149w5150w(0) <= NOT wire_y_pipeff_6_w_q_range5149w(0);
	wire_y_pipeff_6_w_lg_w_q_range5155w5156w(0) <= NOT wire_y_pipeff_6_w_q_range5155w(0);
	wire_y_pipeff_6_w_lg_w_q_range5161w5162w(0) <= NOT wire_y_pipeff_6_w_q_range5161w(0);
	wire_y_pipeff_6_w_lg_w_q_range5167w5168w(0) <= NOT wire_y_pipeff_6_w_q_range5167w(0);
	wire_y_pipeff_6_w_lg_w_q_range5173w5174w(0) <= NOT wire_y_pipeff_6_w_q_range5173w(0);
	wire_y_pipeff_6_w_lg_w_q_range5179w5180w(0) <= NOT wire_y_pipeff_6_w_q_range5179w(0);
	wire_y_pipeff_6_w_lg_w_q_range5185w5186w(0) <= NOT wire_y_pipeff_6_w_q_range5185w(0);
	wire_y_pipeff_6_w_lg_w_q_range5191w5192w(0) <= NOT wire_y_pipeff_6_w_q_range5191w(0);
	wire_y_pipeff_6_w_lg_w_q_range5197w5198w(0) <= NOT wire_y_pipeff_6_w_q_range5197w(0);
	wire_y_pipeff_6_w_lg_w_q_range5203w5204w(0) <= NOT wire_y_pipeff_6_w_q_range5203w(0);
	wire_y_pipeff_6_w_lg_w_q_range5209w5210w(0) <= NOT wire_y_pipeff_6_w_q_range5209w(0);
	wire_y_pipeff_6_w_lg_w_q_range5215w5216w(0) <= NOT wire_y_pipeff_6_w_q_range5215w(0);
	wire_y_pipeff_6_w_lg_w_q_range5221w5222w(0) <= NOT wire_y_pipeff_6_w_q_range5221w(0);
	wire_y_pipeff_6_w_lg_w_q_range5227w5228w(0) <= NOT wire_y_pipeff_6_w_q_range5227w(0);
	wire_y_pipeff_6_w_lg_w_q_range5233w5234w(0) <= NOT wire_y_pipeff_6_w_q_range5233w(0);
	wire_y_pipeff_6_w_lg_w_q_range5239w5240w(0) <= NOT wire_y_pipeff_6_w_q_range5239w(0);
	wire_y_pipeff_6_w_lg_w_q_range5245w5246w(0) <= NOT wire_y_pipeff_6_w_q_range5245w(0);
	wire_y_pipeff_6_w_lg_w_q_range5055w5056w(0) <= NOT wire_y_pipeff_6_w_q_range5055w(0);
	wire_y_pipeff_6_w_lg_w_q_range5090w5091w(0) <= NOT wire_y_pipeff_6_w_q_range5090w(0);
	wire_y_pipeff_6_w_lg_w_q_range5095w5096w(0) <= NOT wire_y_pipeff_6_w_q_range5095w(0);
	wire_y_pipeff_6_w_lg_w_q_range5101w5102w(0) <= NOT wire_y_pipeff_6_w_q_range5101w(0);
	wire_y_pipeff_6_w_lg_w_q_range5107w5108w(0) <= NOT wire_y_pipeff_6_w_q_range5107w(0);
	wire_y_pipeff_6_w_q_range5113w(0) <= y_pipeff_6(10);
	wire_y_pipeff_6_w_q_range5119w(0) <= y_pipeff_6(11);
	wire_y_pipeff_6_w_q_range5125w(0) <= y_pipeff_6(12);
	wire_y_pipeff_6_w_q_range5131w(0) <= y_pipeff_6(13);
	wire_y_pipeff_6_w_q_range5137w(0) <= y_pipeff_6(14);
	wire_y_pipeff_6_w_q_range5143w(0) <= y_pipeff_6(15);
	wire_y_pipeff_6_w_q_range5149w(0) <= y_pipeff_6(16);
	wire_y_pipeff_6_w_q_range5155w(0) <= y_pipeff_6(17);
	wire_y_pipeff_6_w_q_range5161w(0) <= y_pipeff_6(18);
	wire_y_pipeff_6_w_q_range5167w(0) <= y_pipeff_6(19);
	wire_y_pipeff_6_w_q_range5173w(0) <= y_pipeff_6(20);
	wire_y_pipeff_6_w_q_range5179w(0) <= y_pipeff_6(21);
	wire_y_pipeff_6_w_q_range5185w(0) <= y_pipeff_6(22);
	wire_y_pipeff_6_w_q_range5191w(0) <= y_pipeff_6(23);
	wire_y_pipeff_6_w_q_range5197w(0) <= y_pipeff_6(24);
	wire_y_pipeff_6_w_q_range5203w(0) <= y_pipeff_6(25);
	wire_y_pipeff_6_w_q_range5209w(0) <= y_pipeff_6(26);
	wire_y_pipeff_6_w_q_range5215w(0) <= y_pipeff_6(27);
	wire_y_pipeff_6_w_q_range5221w(0) <= y_pipeff_6(28);
	wire_y_pipeff_6_w_q_range5227w(0) <= y_pipeff_6(29);
	wire_y_pipeff_6_w_q_range5233w(0) <= y_pipeff_6(30);
	wire_y_pipeff_6_w_q_range5239w(0) <= y_pipeff_6(31);
	wire_y_pipeff_6_w_q_range5245w(0) <= y_pipeff_6(32);
	wire_y_pipeff_6_w_q_range5055w(0) <= y_pipeff_6(33);
	wire_y_pipeff_6_w_q_range5090w(0) <= y_pipeff_6(6);
	wire_y_pipeff_6_w_q_range5095w(0) <= y_pipeff_6(7);
	wire_y_pipeff_6_w_q_range5101w(0) <= y_pipeff_6(8);
	wire_y_pipeff_6_w_q_range5107w(0) <= y_pipeff_6(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_7 <= y_pipenode_7_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_7_w_lg_w_q_range5938w5939w(0) <= NOT wire_y_pipeff_7_w_q_range5938w(0);
	wire_y_pipeff_7_w_lg_w_q_range5944w5945w(0) <= NOT wire_y_pipeff_7_w_q_range5944w(0);
	wire_y_pipeff_7_w_lg_w_q_range5950w5951w(0) <= NOT wire_y_pipeff_7_w_q_range5950w(0);
	wire_y_pipeff_7_w_lg_w_q_range5956w5957w(0) <= NOT wire_y_pipeff_7_w_q_range5956w(0);
	wire_y_pipeff_7_w_lg_w_q_range5962w5963w(0) <= NOT wire_y_pipeff_7_w_q_range5962w(0);
	wire_y_pipeff_7_w_lg_w_q_range5968w5969w(0) <= NOT wire_y_pipeff_7_w_q_range5968w(0);
	wire_y_pipeff_7_w_lg_w_q_range5974w5975w(0) <= NOT wire_y_pipeff_7_w_q_range5974w(0);
	wire_y_pipeff_7_w_lg_w_q_range5980w5981w(0) <= NOT wire_y_pipeff_7_w_q_range5980w(0);
	wire_y_pipeff_7_w_lg_w_q_range5986w5987w(0) <= NOT wire_y_pipeff_7_w_q_range5986w(0);
	wire_y_pipeff_7_w_lg_w_q_range5992w5993w(0) <= NOT wire_y_pipeff_7_w_q_range5992w(0);
	wire_y_pipeff_7_w_lg_w_q_range5998w5999w(0) <= NOT wire_y_pipeff_7_w_q_range5998w(0);
	wire_y_pipeff_7_w_lg_w_q_range6004w6005w(0) <= NOT wire_y_pipeff_7_w_q_range6004w(0);
	wire_y_pipeff_7_w_lg_w_q_range6010w6011w(0) <= NOT wire_y_pipeff_7_w_q_range6010w(0);
	wire_y_pipeff_7_w_lg_w_q_range6016w6017w(0) <= NOT wire_y_pipeff_7_w_q_range6016w(0);
	wire_y_pipeff_7_w_lg_w_q_range6022w6023w(0) <= NOT wire_y_pipeff_7_w_q_range6022w(0);
	wire_y_pipeff_7_w_lg_w_q_range6028w6029w(0) <= NOT wire_y_pipeff_7_w_q_range6028w(0);
	wire_y_pipeff_7_w_lg_w_q_range6034w6035w(0) <= NOT wire_y_pipeff_7_w_q_range6034w(0);
	wire_y_pipeff_7_w_lg_w_q_range6040w6041w(0) <= NOT wire_y_pipeff_7_w_q_range6040w(0);
	wire_y_pipeff_7_w_lg_w_q_range6046w6047w(0) <= NOT wire_y_pipeff_7_w_q_range6046w(0);
	wire_y_pipeff_7_w_lg_w_q_range6052w6053w(0) <= NOT wire_y_pipeff_7_w_q_range6052w(0);
	wire_y_pipeff_7_w_lg_w_q_range6058w6059w(0) <= NOT wire_y_pipeff_7_w_q_range6058w(0);
	wire_y_pipeff_7_w_lg_w_q_range6064w6065w(0) <= NOT wire_y_pipeff_7_w_q_range6064w(0);
	wire_y_pipeff_7_w_lg_w_q_range6070w6071w(0) <= NOT wire_y_pipeff_7_w_q_range6070w(0);
	wire_y_pipeff_7_w_lg_w_q_range5882w5883w(0) <= NOT wire_y_pipeff_7_w_q_range5882w(0);
	wire_y_pipeff_7_w_lg_w_q_range5921w5922w(0) <= NOT wire_y_pipeff_7_w_q_range5921w(0);
	wire_y_pipeff_7_w_lg_w_q_range5926w5927w(0) <= NOT wire_y_pipeff_7_w_q_range5926w(0);
	wire_y_pipeff_7_w_lg_w_q_range5932w5933w(0) <= NOT wire_y_pipeff_7_w_q_range5932w(0);
	wire_y_pipeff_7_w_q_range5938w(0) <= y_pipeff_7(10);
	wire_y_pipeff_7_w_q_range5944w(0) <= y_pipeff_7(11);
	wire_y_pipeff_7_w_q_range5950w(0) <= y_pipeff_7(12);
	wire_y_pipeff_7_w_q_range5956w(0) <= y_pipeff_7(13);
	wire_y_pipeff_7_w_q_range5962w(0) <= y_pipeff_7(14);
	wire_y_pipeff_7_w_q_range5968w(0) <= y_pipeff_7(15);
	wire_y_pipeff_7_w_q_range5974w(0) <= y_pipeff_7(16);
	wire_y_pipeff_7_w_q_range5980w(0) <= y_pipeff_7(17);
	wire_y_pipeff_7_w_q_range5986w(0) <= y_pipeff_7(18);
	wire_y_pipeff_7_w_q_range5992w(0) <= y_pipeff_7(19);
	wire_y_pipeff_7_w_q_range5998w(0) <= y_pipeff_7(20);
	wire_y_pipeff_7_w_q_range6004w(0) <= y_pipeff_7(21);
	wire_y_pipeff_7_w_q_range6010w(0) <= y_pipeff_7(22);
	wire_y_pipeff_7_w_q_range6016w(0) <= y_pipeff_7(23);
	wire_y_pipeff_7_w_q_range6022w(0) <= y_pipeff_7(24);
	wire_y_pipeff_7_w_q_range6028w(0) <= y_pipeff_7(25);
	wire_y_pipeff_7_w_q_range6034w(0) <= y_pipeff_7(26);
	wire_y_pipeff_7_w_q_range6040w(0) <= y_pipeff_7(27);
	wire_y_pipeff_7_w_q_range6046w(0) <= y_pipeff_7(28);
	wire_y_pipeff_7_w_q_range6052w(0) <= y_pipeff_7(29);
	wire_y_pipeff_7_w_q_range6058w(0) <= y_pipeff_7(30);
	wire_y_pipeff_7_w_q_range6064w(0) <= y_pipeff_7(31);
	wire_y_pipeff_7_w_q_range6070w(0) <= y_pipeff_7(32);
	wire_y_pipeff_7_w_q_range5882w(0) <= y_pipeff_7(33);
	wire_y_pipeff_7_w_q_range5921w(0) <= y_pipeff_7(7);
	wire_y_pipeff_7_w_q_range5926w(0) <= y_pipeff_7(8);
	wire_y_pipeff_7_w_q_range5932w(0) <= y_pipeff_7(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_8 <= y_pipenode_8_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_8_w_lg_w_q_range6758w6759w(0) <= NOT wire_y_pipeff_8_w_q_range6758w(0);
	wire_y_pipeff_8_w_lg_w_q_range6764w6765w(0) <= NOT wire_y_pipeff_8_w_q_range6764w(0);
	wire_y_pipeff_8_w_lg_w_q_range6770w6771w(0) <= NOT wire_y_pipeff_8_w_q_range6770w(0);
	wire_y_pipeff_8_w_lg_w_q_range6776w6777w(0) <= NOT wire_y_pipeff_8_w_q_range6776w(0);
	wire_y_pipeff_8_w_lg_w_q_range6782w6783w(0) <= NOT wire_y_pipeff_8_w_q_range6782w(0);
	wire_y_pipeff_8_w_lg_w_q_range6788w6789w(0) <= NOT wire_y_pipeff_8_w_q_range6788w(0);
	wire_y_pipeff_8_w_lg_w_q_range6794w6795w(0) <= NOT wire_y_pipeff_8_w_q_range6794w(0);
	wire_y_pipeff_8_w_lg_w_q_range6800w6801w(0) <= NOT wire_y_pipeff_8_w_q_range6800w(0);
	wire_y_pipeff_8_w_lg_w_q_range6806w6807w(0) <= NOT wire_y_pipeff_8_w_q_range6806w(0);
	wire_y_pipeff_8_w_lg_w_q_range6812w6813w(0) <= NOT wire_y_pipeff_8_w_q_range6812w(0);
	wire_y_pipeff_8_w_lg_w_q_range6818w6819w(0) <= NOT wire_y_pipeff_8_w_q_range6818w(0);
	wire_y_pipeff_8_w_lg_w_q_range6824w6825w(0) <= NOT wire_y_pipeff_8_w_q_range6824w(0);
	wire_y_pipeff_8_w_lg_w_q_range6830w6831w(0) <= NOT wire_y_pipeff_8_w_q_range6830w(0);
	wire_y_pipeff_8_w_lg_w_q_range6836w6837w(0) <= NOT wire_y_pipeff_8_w_q_range6836w(0);
	wire_y_pipeff_8_w_lg_w_q_range6842w6843w(0) <= NOT wire_y_pipeff_8_w_q_range6842w(0);
	wire_y_pipeff_8_w_lg_w_q_range6848w6849w(0) <= NOT wire_y_pipeff_8_w_q_range6848w(0);
	wire_y_pipeff_8_w_lg_w_q_range6854w6855w(0) <= NOT wire_y_pipeff_8_w_q_range6854w(0);
	wire_y_pipeff_8_w_lg_w_q_range6860w6861w(0) <= NOT wire_y_pipeff_8_w_q_range6860w(0);
	wire_y_pipeff_8_w_lg_w_q_range6866w6867w(0) <= NOT wire_y_pipeff_8_w_q_range6866w(0);
	wire_y_pipeff_8_w_lg_w_q_range6872w6873w(0) <= NOT wire_y_pipeff_8_w_q_range6872w(0);
	wire_y_pipeff_8_w_lg_w_q_range6878w6879w(0) <= NOT wire_y_pipeff_8_w_q_range6878w(0);
	wire_y_pipeff_8_w_lg_w_q_range6884w6885w(0) <= NOT wire_y_pipeff_8_w_q_range6884w(0);
	wire_y_pipeff_8_w_lg_w_q_range6890w6891w(0) <= NOT wire_y_pipeff_8_w_q_range6890w(0);
	wire_y_pipeff_8_w_lg_w_q_range6704w6705w(0) <= NOT wire_y_pipeff_8_w_q_range6704w(0);
	wire_y_pipeff_8_w_lg_w_q_range6747w6748w(0) <= NOT wire_y_pipeff_8_w_q_range6747w(0);
	wire_y_pipeff_8_w_lg_w_q_range6752w6753w(0) <= NOT wire_y_pipeff_8_w_q_range6752w(0);
	wire_y_pipeff_8_w_q_range6758w(0) <= y_pipeff_8(10);
	wire_y_pipeff_8_w_q_range6764w(0) <= y_pipeff_8(11);
	wire_y_pipeff_8_w_q_range6770w(0) <= y_pipeff_8(12);
	wire_y_pipeff_8_w_q_range6776w(0) <= y_pipeff_8(13);
	wire_y_pipeff_8_w_q_range6782w(0) <= y_pipeff_8(14);
	wire_y_pipeff_8_w_q_range6788w(0) <= y_pipeff_8(15);
	wire_y_pipeff_8_w_q_range6794w(0) <= y_pipeff_8(16);
	wire_y_pipeff_8_w_q_range6800w(0) <= y_pipeff_8(17);
	wire_y_pipeff_8_w_q_range6806w(0) <= y_pipeff_8(18);
	wire_y_pipeff_8_w_q_range6812w(0) <= y_pipeff_8(19);
	wire_y_pipeff_8_w_q_range6818w(0) <= y_pipeff_8(20);
	wire_y_pipeff_8_w_q_range6824w(0) <= y_pipeff_8(21);
	wire_y_pipeff_8_w_q_range6830w(0) <= y_pipeff_8(22);
	wire_y_pipeff_8_w_q_range6836w(0) <= y_pipeff_8(23);
	wire_y_pipeff_8_w_q_range6842w(0) <= y_pipeff_8(24);
	wire_y_pipeff_8_w_q_range6848w(0) <= y_pipeff_8(25);
	wire_y_pipeff_8_w_q_range6854w(0) <= y_pipeff_8(26);
	wire_y_pipeff_8_w_q_range6860w(0) <= y_pipeff_8(27);
	wire_y_pipeff_8_w_q_range6866w(0) <= y_pipeff_8(28);
	wire_y_pipeff_8_w_q_range6872w(0) <= y_pipeff_8(29);
	wire_y_pipeff_8_w_q_range6878w(0) <= y_pipeff_8(30);
	wire_y_pipeff_8_w_q_range6884w(0) <= y_pipeff_8(31);
	wire_y_pipeff_8_w_q_range6890w(0) <= y_pipeff_8(32);
	wire_y_pipeff_8_w_q_range6704w(0) <= y_pipeff_8(33);
	wire_y_pipeff_8_w_q_range6747w(0) <= y_pipeff_8(8);
	wire_y_pipeff_8_w_q_range6752w(0) <= y_pipeff_8(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_9 <= y_pipenode_9_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_9_w_lg_w_q_range7573w7574w(0) <= NOT wire_y_pipeff_9_w_q_range7573w(0);
	wire_y_pipeff_9_w_lg_w_q_range7579w7580w(0) <= NOT wire_y_pipeff_9_w_q_range7579w(0);
	wire_y_pipeff_9_w_lg_w_q_range7585w7586w(0) <= NOT wire_y_pipeff_9_w_q_range7585w(0);
	wire_y_pipeff_9_w_lg_w_q_range7591w7592w(0) <= NOT wire_y_pipeff_9_w_q_range7591w(0);
	wire_y_pipeff_9_w_lg_w_q_range7597w7598w(0) <= NOT wire_y_pipeff_9_w_q_range7597w(0);
	wire_y_pipeff_9_w_lg_w_q_range7603w7604w(0) <= NOT wire_y_pipeff_9_w_q_range7603w(0);
	wire_y_pipeff_9_w_lg_w_q_range7609w7610w(0) <= NOT wire_y_pipeff_9_w_q_range7609w(0);
	wire_y_pipeff_9_w_lg_w_q_range7615w7616w(0) <= NOT wire_y_pipeff_9_w_q_range7615w(0);
	wire_y_pipeff_9_w_lg_w_q_range7621w7622w(0) <= NOT wire_y_pipeff_9_w_q_range7621w(0);
	wire_y_pipeff_9_w_lg_w_q_range7627w7628w(0) <= NOT wire_y_pipeff_9_w_q_range7627w(0);
	wire_y_pipeff_9_w_lg_w_q_range7633w7634w(0) <= NOT wire_y_pipeff_9_w_q_range7633w(0);
	wire_y_pipeff_9_w_lg_w_q_range7639w7640w(0) <= NOT wire_y_pipeff_9_w_q_range7639w(0);
	wire_y_pipeff_9_w_lg_w_q_range7645w7646w(0) <= NOT wire_y_pipeff_9_w_q_range7645w(0);
	wire_y_pipeff_9_w_lg_w_q_range7651w7652w(0) <= NOT wire_y_pipeff_9_w_q_range7651w(0);
	wire_y_pipeff_9_w_lg_w_q_range7657w7658w(0) <= NOT wire_y_pipeff_9_w_q_range7657w(0);
	wire_y_pipeff_9_w_lg_w_q_range7663w7664w(0) <= NOT wire_y_pipeff_9_w_q_range7663w(0);
	wire_y_pipeff_9_w_lg_w_q_range7669w7670w(0) <= NOT wire_y_pipeff_9_w_q_range7669w(0);
	wire_y_pipeff_9_w_lg_w_q_range7675w7676w(0) <= NOT wire_y_pipeff_9_w_q_range7675w(0);
	wire_y_pipeff_9_w_lg_w_q_range7681w7682w(0) <= NOT wire_y_pipeff_9_w_q_range7681w(0);
	wire_y_pipeff_9_w_lg_w_q_range7687w7688w(0) <= NOT wire_y_pipeff_9_w_q_range7687w(0);
	wire_y_pipeff_9_w_lg_w_q_range7693w7694w(0) <= NOT wire_y_pipeff_9_w_q_range7693w(0);
	wire_y_pipeff_9_w_lg_w_q_range7699w7700w(0) <= NOT wire_y_pipeff_9_w_q_range7699w(0);
	wire_y_pipeff_9_w_lg_w_q_range7705w7706w(0) <= NOT wire_y_pipeff_9_w_q_range7705w(0);
	wire_y_pipeff_9_w_lg_w_q_range7521w7522w(0) <= NOT wire_y_pipeff_9_w_q_range7521w(0);
	wire_y_pipeff_9_w_lg_w_q_range7568w7569w(0) <= NOT wire_y_pipeff_9_w_q_range7568w(0);
	wire_y_pipeff_9_w_q_range7573w(0) <= y_pipeff_9(10);
	wire_y_pipeff_9_w_q_range7579w(0) <= y_pipeff_9(11);
	wire_y_pipeff_9_w_q_range7585w(0) <= y_pipeff_9(12);
	wire_y_pipeff_9_w_q_range7591w(0) <= y_pipeff_9(13);
	wire_y_pipeff_9_w_q_range7597w(0) <= y_pipeff_9(14);
	wire_y_pipeff_9_w_q_range7603w(0) <= y_pipeff_9(15);
	wire_y_pipeff_9_w_q_range7609w(0) <= y_pipeff_9(16);
	wire_y_pipeff_9_w_q_range7615w(0) <= y_pipeff_9(17);
	wire_y_pipeff_9_w_q_range7621w(0) <= y_pipeff_9(18);
	wire_y_pipeff_9_w_q_range7627w(0) <= y_pipeff_9(19);
	wire_y_pipeff_9_w_q_range7633w(0) <= y_pipeff_9(20);
	wire_y_pipeff_9_w_q_range7639w(0) <= y_pipeff_9(21);
	wire_y_pipeff_9_w_q_range7645w(0) <= y_pipeff_9(22);
	wire_y_pipeff_9_w_q_range7651w(0) <= y_pipeff_9(23);
	wire_y_pipeff_9_w_q_range7657w(0) <= y_pipeff_9(24);
	wire_y_pipeff_9_w_q_range7663w(0) <= y_pipeff_9(25);
	wire_y_pipeff_9_w_q_range7669w(0) <= y_pipeff_9(26);
	wire_y_pipeff_9_w_q_range7675w(0) <= y_pipeff_9(27);
	wire_y_pipeff_9_w_q_range7681w(0) <= y_pipeff_9(28);
	wire_y_pipeff_9_w_q_range7687w(0) <= y_pipeff_9(29);
	wire_y_pipeff_9_w_q_range7693w(0) <= y_pipeff_9(30);
	wire_y_pipeff_9_w_q_range7699w(0) <= y_pipeff_9(31);
	wire_y_pipeff_9_w_q_range7705w(0) <= y_pipeff_9(32);
	wire_y_pipeff_9_w_q_range7521w(0) <= y_pipeff_9(33);
	wire_y_pipeff_9_w_q_range7568w(0) <= y_pipeff_9(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_0 <= radians_load_node_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_1 <= wire_z_pipeff1_sub_result;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_1_w_q_range1421w(0) <= z_pipeff_1(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_10 <= z_pipenode_10_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_10_w_q_range8864w(0) <= z_pipeff_10(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_11 <= z_pipenode_11_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_11_w_q_range9666w(0) <= z_pipeff_11(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_12 <= z_pipenode_12_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_12_w_q_range10463w(0) <= z_pipeff_12(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_13 <= z_pipenode_13_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_2 <= z_pipenode_2_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_2_w_q_range2268w(0) <= z_pipeff_2(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_3 <= z_pipenode_3_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_3_w_q_range3110w(0) <= z_pipeff_3(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_4 <= z_pipenode_4_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_4_w_q_range3947w(0) <= z_pipeff_4(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_5 <= z_pipenode_5_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_5_w_q_range4779w(0) <= z_pipeff_5(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_6 <= z_pipenode_6_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_6_w_q_range5606w(0) <= z_pipeff_6(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_7 <= z_pipenode_7_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_7_w_q_range6428w(0) <= z_pipeff_7(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_8 <= z_pipenode_8_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_8_w_q_range7245w(0) <= z_pipeff_8(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_9 <= z_pipenode_9_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_9_w_q_range8057w(0) <= z_pipeff_9(33);
	wire_sincos_add_cin <= wire_sincosbitff_w_lg_w_q_range10746w10747w(0);
	sincos_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => wire_sincos_add_cin,
		dataa => delay_pipe_w,
		datab => post_estimate_w,
		result => wire_sincos_add_result
	  );
	x_pipenode_10_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_9(33),
		dataa => x_pipeff_9,
		datab => x_subnode_10_w,
		result => wire_x_pipenode_10_add_result
	  );
	x_pipenode_11_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_10(33),
		dataa => x_pipeff_10,
		datab => x_subnode_11_w,
		result => wire_x_pipenode_11_add_result
	  );
	x_pipenode_12_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_11(33),
		dataa => x_pipeff_11,
		datab => x_subnode_12_w,
		result => wire_x_pipenode_12_add_result
	  );
	x_pipenode_13_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_12(33),
		dataa => x_pipeff_12,
		datab => x_subnode_13_w,
		result => wire_x_pipenode_13_add_result
	  );
	x_pipenode_2_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_1(33),
		dataa => x_pipeff_1,
		datab => x_subnode_2_w,
		result => wire_x_pipenode_2_add_result
	  );
	x_pipenode_3_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_2(33),
		dataa => x_pipeff_2,
		datab => x_subnode_3_w,
		result => wire_x_pipenode_3_add_result
	  );
	x_pipenode_4_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_3(33),
		dataa => x_pipeff_3,
		datab => x_subnode_4_w,
		result => wire_x_pipenode_4_add_result
	  );
	x_pipenode_5_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_4(33),
		dataa => x_pipeff_4,
		datab => x_subnode_5_w,
		result => wire_x_pipenode_5_add_result
	  );
	x_pipenode_6_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_5(33),
		dataa => x_pipeff_5,
		datab => x_subnode_6_w,
		result => wire_x_pipenode_6_add_result
	  );
	x_pipenode_7_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_6(33),
		dataa => x_pipeff_6,
		datab => x_subnode_7_w,
		result => wire_x_pipenode_7_add_result
	  );
	x_pipenode_8_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_7(33),
		dataa => x_pipeff_7,
		datab => x_subnode_8_w,
		result => wire_x_pipenode_8_add_result
	  );
	x_pipenode_9_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_8(33),
		dataa => x_pipeff_8,
		datab => x_subnode_9_w,
		result => wire_x_pipenode_9_add_result
	  );
	y_pipeff1_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		dataa => y_pipeff_0,
		datab => y_subnode_1_w,
		result => wire_y_pipeff1_add_result
	  );
	y_pipenode_10_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_9(33),
		dataa => y_pipeff_9,
		datab => y_subnode_10_w,
		result => wire_y_pipenode_10_add_result
	  );
	y_pipenode_11_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_10(33),
		dataa => y_pipeff_10,
		datab => y_subnode_11_w,
		result => wire_y_pipenode_11_add_result
	  );
	y_pipenode_12_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_11(33),
		dataa => y_pipeff_11,
		datab => y_subnode_12_w,
		result => wire_y_pipenode_12_add_result
	  );
	y_pipenode_13_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_12(33),
		dataa => y_pipeff_12,
		datab => y_subnode_13_w,
		result => wire_y_pipenode_13_add_result
	  );
	y_pipenode_2_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_1(33),
		dataa => y_pipeff_1,
		datab => y_subnode_2_w,
		result => wire_y_pipenode_2_add_result
	  );
	y_pipenode_3_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_2(33),
		dataa => y_pipeff_2,
		datab => y_subnode_3_w,
		result => wire_y_pipenode_3_add_result
	  );
	y_pipenode_4_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_3(33),
		dataa => y_pipeff_3,
		datab => y_subnode_4_w,
		result => wire_y_pipenode_4_add_result
	  );
	y_pipenode_5_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_4(33),
		dataa => y_pipeff_4,
		datab => y_subnode_5_w,
		result => wire_y_pipenode_5_add_result
	  );
	y_pipenode_6_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_5(33),
		dataa => y_pipeff_5,
		datab => y_subnode_6_w,
		result => wire_y_pipenode_6_add_result
	  );
	y_pipenode_7_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_6(33),
		dataa => y_pipeff_6,
		datab => y_subnode_7_w,
		result => wire_y_pipenode_7_add_result
	  );
	y_pipenode_8_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_7(33),
		dataa => y_pipeff_7,
		datab => y_subnode_8_w,
		result => wire_y_pipenode_8_add_result
	  );
	y_pipenode_9_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_8(33),
		dataa => y_pipeff_8,
		datab => y_subnode_9_w,
		result => wire_y_pipenode_9_add_result
	  );
	z_pipeff1_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		dataa => z_pipeff_0,
		datab => atannode_0_w,
		result => wire_z_pipeff1_sub_result
	  );
	z_pipenode_10_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_9(33),
		dataa => z_pipeff_9,
		datab => z_subnode_10_w,
		result => wire_z_pipenode_10_add_result
	  );
	z_pipenode_11_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_10(33),
		dataa => z_pipeff_10,
		datab => z_subnode_11_w,
		result => wire_z_pipenode_11_add_result
	  );
	z_pipenode_12_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_11(33),
		dataa => z_pipeff_11,
		datab => z_subnode_12_w,
		result => wire_z_pipenode_12_add_result
	  );
	z_pipenode_13_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_12(33),
		dataa => z_pipeff_12,
		datab => z_subnode_13_w,
		result => wire_z_pipenode_13_add_result
	  );
	z_pipenode_2_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_1(33),
		dataa => z_pipeff_1,
		datab => z_subnode_2_w,
		result => wire_z_pipenode_2_add_result
	  );
	z_pipenode_3_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_2(33),
		dataa => z_pipeff_2,
		datab => z_subnode_3_w,
		result => wire_z_pipenode_3_add_result
	  );
	z_pipenode_4_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_3(33),
		dataa => z_pipeff_3,
		datab => z_subnode_4_w,
		result => wire_z_pipenode_4_add_result
	  );
	z_pipenode_5_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_4(33),
		dataa => z_pipeff_4,
		datab => z_subnode_5_w,
		result => wire_z_pipenode_5_add_result
	  );
	z_pipenode_6_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_5(33),
		dataa => z_pipeff_5,
		datab => z_subnode_6_w,
		result => wire_z_pipenode_6_add_result
	  );
	z_pipenode_7_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_6(33),
		dataa => z_pipeff_6,
		datab => z_subnode_7_w,
		result => wire_z_pipenode_7_add_result
	  );
	z_pipenode_8_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_7(33),
		dataa => z_pipeff_7,
		datab => z_subnode_8_w,
		result => wire_z_pipenode_8_add_result
	  );
	z_pipenode_9_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		cin => z_pipeff_8(33),
		dataa => z_pipeff_8,
		datab => z_subnode_9_w,
		result => wire_z_pipenode_9_add_result
	  );
	cmx :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTHA => 34,
		LPM_WIDTHB => 34,
		LPM_WIDTHP => 68
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => multiplier_input_w,
		datab => z_pipeff_13,
		result => wire_cmx_result
	  );

 END RTL; --sinhw_altfp_sincos_cordic_m_e5e


--altfp_sincos_range CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" WIDTH_EXP=8 WIDTH_MAN=23 aclr circle clken clock data negcircle
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END


--altfp_sincos_srrt CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" address basefraction incexponent incmantissa
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_mux 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_srrt_koa IS 
	 PORT 
	 ( 
		 address	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 basefraction	:	OUT  STD_LOGIC_VECTOR (35 DOWNTO 0);
		 incexponent	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 incmantissa	:	OUT  STD_LOGIC_VECTOR (55 DOWNTO 0)
	 ); 
 END sinhw_altfp_sincos_srrt_koa;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_srrt_koa IS

	 SIGNAL  wire_mux2_data	:	STD_LOGIC_VECTOR (25599 DOWNTO 0);
	 SIGNAL  wire_mux2_data_2d	:	STD_LOGIC_2D(255 DOWNTO 0, 99 DOWNTO 0);
	 SIGNAL  wire_mux2_result	:	STD_LOGIC_VECTOR (99 DOWNTO 0);
 BEGIN

	basefraction <= wire_mux2_result(35 DOWNTO 0);
	incexponent <= wire_mux2_result(99 DOWNTO 92);
	incmantissa <= wire_mux2_result(91 DOWNTO 36);
	wire_mux2_data <= ( "00000000" & "10011010011011101110000001101101101100010100101011001000" & "00110110" & "1101100010100101011001100101" & "00000001" & "10011010011011101110000001101101101100010100101011010000" & "00011011" & "0110110001010010101100110010" & "00000000" & "10100110100110111011100000011011011011000101001010111000" & "00001101" & "1011011000101001010110011001" & "00000001" & "10100110100110111011100000011011011011000101001010110000" & "00000110" & "1101101100010100101011001101" & "00000000" & "10101001101001101110111000000110110110110001010010110000" & "00000011" & "0110110110001010010101100110" & "00000000" & "11010100110100110111011100000011011011011000101001100000" & "10000001" & "1011011011000101001010110011" & "00000000" & "11101010011010011011101110000001101101101100010100011000" & "11000000" & "1101101101100010100101011010" & "00000000" & "11110101001101001101110111000000110110110110001010011000" & "11100000" & "0110110110110001010010101101" & "00000000" & "11111010100110100110111011100000011011011011000101010000" & "01110000" & "0011011011011000101001010110" & "00000001" & "11111010100110100110111011100000011011011011000101010000" & "10111000" & "0001101101101100010100101011" & "00000010" & "11111010100110100110111011100000011011011011000101010000" & "11011100" & "0000110110110110001010010110" & "00000011" & "11111010100110100110111011100000011011011011000100101000" & "11101110" & "0000011011011011000101001011" & "00000000" & "10001111101010011010011011101110000001101101101100011000" & "01110111" & "0000001101101101100010100101" & "00000001" & "10001111101010011010011011101110000001101101101100100000" & "10111011" & "1000000110110110110001010011" & "00000000" & "10100011111010100110100110111011100000011011011011001000" & "11011101" & "1100000011011011011000101001" & "00000000" & "11010001111101010011010011011101110000001101101101010000" & "01101110" & "1110000001101101101100010101" & "00000000" & "11101000111110101001101001101110111000000110110110111000" & "00110111" & "0111000000110110110110001010"
 & "00000000" & "11110100011111010100110100110111011100000011011011011000" & "10011011" & "1011100000011011011011000101" & "00000000" & "11111010001111101010011010011011101110000001101101101000" & "01001101" & "1101110000001101101101100011" & "00000001" & "11111010001111101010011010011011101110000001101110000000" & "10100110" & "1110111000000110110110110001" & "00000000" & "10111110100011111010100110100110111011100000011011100000" & "11010011" & "0111011100000011011011011001" & "00000001" & "10111110100011111010100110100110111011100000011011101000" & "01101001" & "1011101110000001101101101100" & "00000000" & "10101111101000111110101001101001101110111000000110111000" & "00110100" & "1101110111000000110110110110" & "00000001" & "10101111101000111110101001101001101110111000000110110000" & "10011010" & "0110111011100000011011011011" & "00000000" & "10101011111010001111101010011010011011101110000001110000" & "01001101" & "0011011101110000001101101110" & "00000000" & "11010101111101000111110101001101001101110111000000111000" & "10100110" & "1001101110111000000110110111" & "00000000" & "11101010111110100011111010100110100110111011100000110000" & "01010011" & "0100110111011100000011011011" & "00000001" & "11101010111110100011111010100110100110111011100000100000" & "10101001" & "1010011011101110000001101110" & "00000010" & "11101010111110100011111010100110100110111011011111111000" & "11010100" & "1101001101110111000000110111" & "00000000" & "10011101010111110100011111010100110100110111011100000000" & "11101010" & "0110100110111011100000011011" & "00000001" & "10011101010111110100011111010100110100110111011100011000" & "11110101" & "0011010011011101110000001110" & "00000010" & "10011101010111110100011111010100110100110111011100011000" & "11111010" & "1001101001101110111000000111" & "00000011" & "10011101010111110100011111010100110100110111011100011000" & "01111101" & "0100110100110111011100000011" & "00000100" & "10011101010111110100011111010100110100110111011110010000" & "00111110" & "1010011010011011101110000010" & "00000000"
 & "10000100111010101111101000111110101001101001101111000000" & "00011111" & "0101001101001101110111000001" & "00000000" & "11000010011101010111110100011111010100110100110111011000" & "10001111" & "1010100110100110111011100000" & "00000000" & "11100001001110101011111010001111101010011010011011110000" & "01000111" & "1101010011010011011101110000" & "00000000" & "11110000100111010101111101000111110101001101001110000000" & "10100011" & "1110101001101001101110111000" & "00000000" & "11111000010011101010111110100011111010100110100110111000" & "11010001" & "1111010100110100110111011100" & "00000000" & "11111100001001110101011111010001111101010011010011011000" & "11101000" & "1111101010011010011011101110" & "00000000" & "11111110000100111010101111101000111110101001101001110000" & "11110100" & "0111110101001101001101110111" & "00000001" & "11111110000100111010101111101000111110101001101010000000" & "11111010" & "0011111010100110100110111100" & "00000010" & "11111110000100111010101111101000111110101001101001110000" & "01111101" & "0001111101010011010011011110" & "00000000" & "10011111110000100111010101111101000111110101001101011000" & "10111110" & "1000111110101001101001101111" & "00000001" & "10011111110000100111010101111101000111110101001101100000" & "01011111" & "0100011111010100110100110111" & "00000000" & "10100111111100001001110101011111010001111101010011010000" & "10101111" & "1010001111101010011010011100" & "00000001" & "10100111111100001001110101011111010001111101010011100000" & "01010111" & "1101000111110101001101001110" & "00000010" & "10100111111100001001110101011111010001111101010011010000" & "10101011" & "1110100011111010100110100111" & "00000000" & "10010100111111100001001110101011111010001111101010011000" & "11010101" & "1111010001111101010011010011" & "00000001" & "10010100111111100001001110101011111010001111101010101000" & "11101010" & "1111101000111110101001101010" & "00000000" & "10100101001111111000010011101010111110100011111010101000" & "01110101" & "0111110100011111010100110101" & "00000001" & "10100101001111111000010011101010111110100011111010101000"
 & "00111010" & "1011111010001111101010011010" & "00000000" & "10101001010011111110000100111010101111101000111110101000" & "10011101" & "0101111101000111110101001101" & "00000001" & "10101001010011111110000100111010101111101000111110111000" & "01001110" & "1010111110100011111010100111" & "00000010" & "10101001010011111110000100111010101111101000111110111000" & "00100111" & "0101011111010001111101010011" & "00000011" & "10101001010011111110000100111010101111101000111110111000" & "00010011" & "1010101111101000111110101010" & "00000100" & "10101001010011111110000100111010101111101000111110111000" & "00001001" & "1101010111110100011111010101" & "00000101" & "10101001010011111110000100111010101111101001000000110000" & "10000100" & "1110101011111010001111101010" & "00000000" & "10000010101001010011111110000100111010101111101001001000" & "11000010" & "0111010101111101000111110101" & "00000001" & "10000010101001010011111110000100111010101111101001010000" & "11100001" & "0011101010111110100011111011" & "00000010" & "10000010101001010011111110000100111010101111101000111000" & "11110000" & "1001110101011111010001111101" & "00000011" & "10000010101001010011111110000100111010101111101001100000" & "11111000" & "0100111010101111101000111111" & "00000000" & "10001000001010100101001111111000010011101010111110100000" & "11111100" & "0010011101010111110100011111" & "00000001" & "10001000001010100101001111111000010011101010111110100000" & "11111110" & "0001001110101011111010010000" & "00000010" & "10001000001010100101001111111000010011101010111110100000" & "01111111" & "0000100111010101111101001000" & "00000000" & "10010001000001010100101001111111000010011101011000010000" & "00111111" & "1000010011101010111110100100" & "00000000" & "11001000100000101010010100111111100001001110101011111000" & "10011111" & "1100001001110101011111010010" & "00000000" & "11100100010000010101001010011111110000100111010101111000" & "01001111" & "1110000100111010101111101001" & "00000001" & "11100100010000010101001010011111110000100111010101110000" & "10100111"
 & "1111000010011101010111110100" & "00000010" & "11100100010000010101001010011111110000100111010110001000" & "01010011" & "1111100001001110101011111010" & "00000000" & "10011100100010000010101001010011111110000100111010111000" & "00101001" & "1111110000100111010101111101" & "00000001" & "10011100100010000010101001010011111110000100111010111000" & "10010100" & "1111111000010011101010111111" & "00000010" & "10011100100010000010101001010011111110000100111010110000" & "01001010" & "0111111100001001110101011111" & "00000000" & "10010011100100010000010101001010011111110000100111011000" & "10100101" & "0011111110000100111010110000" & "00000000" & "11001001110010001000001010100101001111111000010011101000" & "01010010" & "1001111111000010011101011000" & "00000000" & "11100100111001000100000101010010100111111100001001111000" & "10101001" & "0100111111100001001110101100" & "00000001" & "11100100111001000100000101010010100111111100001001101000" & "01010100" & "1010011111110000100111010110" & "00000000" & "10111001001110010001000001010100101001111111000010011000" & "00101010" & "0101001111111000010011101011" & "00000000" & "11011100100111001000100000101010010100111111100001011000" & "00010101" & "0010100111111100001001110101" & "00000001" & "11011100100111001000100000101010010100111111100001011000" & "00001010" & "1001010011111110000100111011" & "00000000" & "10110111001001110010001000001010100101001111111000011000" & "00000101" & "0100101001111111000010011101" & "00000000" & "11011011100100111001000100000101010010100111111100001000" & "10000010" & "1010010100111111100001001111" & "00000001" & "11011011100100111001000100000101010010100111111011111000" & "01000001" & "0101001010011111110000100111" & "00000010" & "11011011100100111001000100000101010010100111111100001000" & "00100000" & "1010100101001111111000010100" & "00000011" & "11011011100100111001000100000101010010100111111100100000" & "00010000" & "0101010010100111111100001010" & "00000100" & "11011011100100111001000100000101010010100111111010111000" & "10001000" & "0010101001010011111110000101"
 & "00000101" & "11011011100100111001000100000101010010100111111001101000" & "01000100" & "0001010100101001111111000010" & "00000000" & "10000011011011100100111001000100000101010010101000000000" & "00100010" & "0000101010010100111111100001" & "00000000" & "11000001101101110010011100100010000010101001010100001000" & "10010001" & "0000010101001010011111110001" & "00000001" & "11000001101101110010011100100010000010101001010011110000" & "11001000" & "1000001010100101001111111000" & "00000010" & "11000001101101110010011100100010000010101001010100001000" & "11100100" & "0100000101010010100111111100" & "00000000" & "10011000001101101110010011100100010000010101001010100000" & "01110010" & "0010000010101001010011111110" & "00000000" & "11001100000110110111001001110010001000001010100101010000" & "00111001" & "0001000001010100101001111111" & "00000000" & "11100110000011011011100100111001000100000101010010101000" & "10011100" & "1000100000101010010101000000" & "00000000" & "11110011000001101101110010011100100010000010101001001000" & "01001110" & "0100010000010101001010100000" & "00000000" & "11111001100000110110111001001110010001000001010100101000" & "00100111" & "0010001000001010100101010000" & "00000001" & "11111001100000110110111001001110010001000001010100101000" & "10010011" & "1001000100000101010010101000" & "00000000" & "10111110011000001101101110010011100100010000010101010000" & "11001001" & "1100100010000010101001010100" & "00000001" & "10111110011000001101101110010011100100010000010101011000" & "11100100" & "1110010001000001010100101010" & "00000010" & "10111110011000001101101110010011100100010000010101000000" & "01110010" & "0111001000100000101010010101" & "00000011" & "10111110011000001101101110010011100100010000010101110000" & "10111001" & "0011100100010000010101001010" & "00000000" & "10001011111001100000110110111001001110010001000001011000" & "11011100" & "1001110010001000001010100101" & "00000001" & "10001011111001100000110110111001001110010001000001010000" & "01101110" & "0100111001000100000101010011" & "00000000"
 & "10100010111110011000001101101110010011100100010000010000" & "10110111" & "0010011100100010000010101001" & "00000001" & "10100010111110011000001101101110010011100100010000011000" & "11011011" & "1001001110010001000001010101" & "00000010" & "10100010111110011000001101101110010011100100010000011000" & "01101101" & "1100100111001000100000101010" & "00000011" & "10100010111110011000001101101110010011100100010000011000" & "00110110" & "1110010011100100010000010101" & "00000100" & "10100010111110011000001101101110010011100100010000011000" & "00011011" & "0111001001110010001000001011" & "00000101" & "10100010111110011000001101101110010011100100010000011000" & "00001101" & "1011100100111001000100000101" & "00000110" & "10100010111110011000001101101110010011100100010000011000" & "00000110" & "1101110010011100100010000011" & "00000111" & "10100010111110011000001101101110010011100100010000011000" & "10000011" & "0110111001001110010001000001" & "00001000" & "10100010111110011000001101101110010011100101100001111000" & "11000001" & "1011011100100111001000100001" & "00001001" & "10100010111110011000001101101110010011100100010000011000" & "01100000" & "1101101110010011100100010000" & "00001010" & "10100010111110011000001101101110010011100100010000011000" & "00110000" & "0110110111001001110010001000" & "00001011" & "10100010111110011000001101101110010011100100010000011000" & "10011000" & "0011011011100100111001000100" & "00001100" & "10100010111110011000001101101110010011100100010000011000" & "11001100" & "0001101101110010011100100010" & "00001101" & "10100010111110011000001101101110010011100100010000011000" & "11100110" & "0000110110111001001110010001" & "00001110" & "10100010111110011000001101101110010011100100010000011000" & "11110011" & "0000011011011100100111001001" & "00001111" & "10100010111110011000001101101110010011100100010000011000" & "11111001" & "1000001101101110010011100100" & "00010000" & "10100010111110011000001101101110010011100100010000011000" & "01111100" & "1100000110110111001001110010" & "00010001" & "10100010111110011000001101101110001001011000010110111000"
 & "10111110" & "0110000011011011100100111001" & "00010010" & "10100010111110011000001101101110010011100100010000011000" & "01011111" & "0011000001101101110010011101" & "00010011" & "10100010111110011000001101101110011000101010001101001000" & "00101111" & "1001100000110110111001001110" & "00010100" & "10100010111110011000001101101110010011100100010000011000" & "00010111" & "1100110000011011011100100111" & "00010101" & "10100010111110011000001101101110010011100100010000011000" & "10001011" & "1110011000001101101110010100" & "00010110" & "10100010111110011000001101101110010011100100010000011000" & "01000101" & "1111001100000110110111001010" & "00010111" & "10100010111110011000001101101110010011100100010000011000" & "10100010" & "1111100110000011011011100101" & "00011000" & "10100010111110011000001101110000110110100010101000101000" & "01010001" & "0111110011000001101101110010" & "00011001" & "10100010111110011000001101101110010011100100010000011000" & "00101000" & "1011111001100000110110111001" & "00011010" & "10100010111110011000001101101110010011100100010000011000" & "00010100" & "0101111100110000011011011101" & "00011011" & "10100010111110011000001101101110010011100100010000011000" & "00001010" & "0010111110011000001101101110" & "00011100" & "10100010111110011000001101101110010011100100010000011000" & "00000101" & "0001011111001100000110110111" & "00011101" & "10100010111110011000001101101110010011100100010000011000" & "00000010" & "1000101111100110000011011100" & "00011110" & "10100010111110011000001101101110010011100100010000011000" & "00000001" & "0100010111110011000001101110" & "00011111" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "1010001011111001100000110111" & "00100000" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0101000101111100110000011011" & "00100001" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0010100010111110011000001110" & "00100010" & "10100010111110011000001101101110010011100100010000011000" & "00000000"
 & "0001010001011111001100000111" & "00100011" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000101000101111100110000011" & "00100100" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000010100010111110011000010" & "00100101" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000001010001011111001100001" & "00100110" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000101000101111100110000" & "00100111" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000010100010111110011000" & "00101000" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000001010001011111001100" & "00101001" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000000101000101111100110" & "00101010" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000000010100010111110011" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
	loop36 : FOR i IN 0 TO 255 GENERATE
		loop37 : FOR j IN 0 TO 99 GENERATE
			wire_mux2_data_2d(i, j) <= wire_mux2_data(i*100+j);
		END GENERATE loop37;
	END GENERATE loop36;
	mux2 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 256,
		LPM_WIDTH => 100,
		LPM_WIDTHS => 8
	  )
	  PORT MAP ( 
		data => wire_mux2_data_2d,
		result => wire_mux2_result,
		sel => address
	  );

 END RTL; --sinhw_altfp_sincos_srrt_koa


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altpriority_encoder_3e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END sinhw_altpriority_encoder_3e8;

 ARCHITECTURE RTL OF sinhw_altpriority_encoder_3e8 IS

 BEGIN

	q(0) <= ( data(1));
	zero <= (NOT (data(0) OR data(1)));

 END RTL; --sinhw_altpriority_encoder_3e8


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altpriority_encoder_3v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END sinhw_altpriority_encoder_3v7;

 ARCHITECTURE RTL OF sinhw_altpriority_encoder_3v7 IS

 BEGIN

	q(0) <= ( data(1));

 END RTL; --sinhw_altpriority_encoder_3v7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altpriority_encoder_6v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END sinhw_altpriority_encoder_6v7;

 ARCHITECTURE RTL OF sinhw_altpriority_encoder_6v7 IS

	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero13017w13018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero13019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero13017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero13019w13020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder9_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  sinhw_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altpriority_encoder_3v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder10_w_lg_zero13017w & wire_altpriority_encoder10_w_lg_w_lg_zero13019w13020w);
	wire_altpriority_encoder10_w_lg_w_lg_zero13017w13018w(0) <= wire_altpriority_encoder10_w_lg_zero13017w(0) AND wire_altpriority_encoder10_q(0);
	wire_altpriority_encoder10_w_lg_zero13019w(0) <= wire_altpriority_encoder10_zero AND wire_altpriority_encoder9_q(0);
	wire_altpriority_encoder10_w_lg_zero13017w(0) <= NOT wire_altpriority_encoder10_zero;
	wire_altpriority_encoder10_w_lg_w_lg_zero13019w13020w(0) <= wire_altpriority_encoder10_w_lg_zero13019w(0) OR wire_altpriority_encoder10_w_lg_w_lg_zero13017w13018w(0);
	altpriority_encoder10 :  sinhw_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder10_q,
		zero => wire_altpriority_encoder10_zero
	  );
	altpriority_encoder9 :  sinhw_altpriority_encoder_3v7
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder9_q
	  );

 END RTL; --sinhw_altpriority_encoder_6v7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altpriority_encoder_6e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END sinhw_altpriority_encoder_6e8;

 ARCHITECTURE RTL OF sinhw_altpriority_encoder_6e8 IS

	 SIGNAL  wire_altpriority_encoder11_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero13035w13036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero13037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero13035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero13037w13038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_zero	:	STD_LOGIC;
	 COMPONENT  sinhw_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder12_w_lg_zero13035w & wire_altpriority_encoder12_w_lg_w_lg_zero13037w13038w);
	zero <= (wire_altpriority_encoder11_zero AND wire_altpriority_encoder12_zero);
	altpriority_encoder11 :  sinhw_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder11_q,
		zero => wire_altpriority_encoder11_zero
	  );
	wire_altpriority_encoder12_w_lg_w_lg_zero13035w13036w(0) <= wire_altpriority_encoder12_w_lg_zero13035w(0) AND wire_altpriority_encoder12_q(0);
	wire_altpriority_encoder12_w_lg_zero13037w(0) <= wire_altpriority_encoder12_zero AND wire_altpriority_encoder11_q(0);
	wire_altpriority_encoder12_w_lg_zero13035w(0) <= NOT wire_altpriority_encoder12_zero;
	wire_altpriority_encoder12_w_lg_w_lg_zero13037w13038w(0) <= wire_altpriority_encoder12_w_lg_zero13037w(0) OR wire_altpriority_encoder12_w_lg_w_lg_zero13035w13036w(0);
	altpriority_encoder12 :  sinhw_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder12_q,
		zero => wire_altpriority_encoder12_zero
	  );

 END RTL; --sinhw_altpriority_encoder_6e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altpriority_encoder_bv7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END sinhw_altpriority_encoder_bv7;

 ARCHITECTURE RTL OF sinhw_altpriority_encoder_bv7 IS

	 SIGNAL  wire_altpriority_encoder7_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_w_lg_zero13008w13009w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_zero13010w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_zero13008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_w_lg_zero13010w13011w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_zero	:	STD_LOGIC;
	 COMPONENT  sinhw_altpriority_encoder_6v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder8_w_lg_zero13008w & wire_altpriority_encoder8_w_lg_w_lg_zero13010w13011w);
	altpriority_encoder7 :  sinhw_altpriority_encoder_6v7
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder7_q
	  );
	loop38 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder8_w_lg_w_lg_zero13008w13009w(i) <= wire_altpriority_encoder8_w_lg_zero13008w(0) AND wire_altpriority_encoder8_q(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder8_w_lg_zero13010w(i) <= wire_altpriority_encoder8_zero AND wire_altpriority_encoder7_q(i);
	END GENERATE loop39;
	wire_altpriority_encoder8_w_lg_zero13008w(0) <= NOT wire_altpriority_encoder8_zero;
	loop40 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder8_w_lg_w_lg_zero13010w13011w(i) <= wire_altpriority_encoder8_w_lg_zero13010w(i) OR wire_altpriority_encoder8_w_lg_w_lg_zero13008w13009w(i);
	END GENERATE loop40;
	altpriority_encoder8 :  sinhw_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder8_q,
		zero => wire_altpriority_encoder8_zero
	  );

 END RTL; --sinhw_altpriority_encoder_bv7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altpriority_encoder_be8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END sinhw_altpriority_encoder_be8;

 ARCHITECTURE RTL OF sinhw_altpriority_encoder_be8 IS

	 SIGNAL  wire_altpriority_encoder13_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero13045w13046w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero13047w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero13045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero13047w13048w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_zero	:	STD_LOGIC;
	 COMPONENT  sinhw_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder14_w_lg_zero13045w & wire_altpriority_encoder14_w_lg_w_lg_zero13047w13048w);
	zero <= (wire_altpriority_encoder13_zero AND wire_altpriority_encoder14_zero);
	altpriority_encoder13 :  sinhw_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder13_q,
		zero => wire_altpriority_encoder13_zero
	  );
	loop41 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero13045w13046w(i) <= wire_altpriority_encoder14_w_lg_zero13045w(0) AND wire_altpriority_encoder14_q(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_zero13047w(i) <= wire_altpriority_encoder14_zero AND wire_altpriority_encoder13_q(i);
	END GENERATE loop42;
	wire_altpriority_encoder14_w_lg_zero13045w(0) <= NOT wire_altpriority_encoder14_zero;
	loop43 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero13047w13048w(i) <= wire_altpriority_encoder14_w_lg_zero13047w(i) OR wire_altpriority_encoder14_w_lg_w_lg_zero13045w13046w(i);
	END GENERATE loop43;
	altpriority_encoder14 :  sinhw_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder14_q,
		zero => wire_altpriority_encoder14_zero
	  );

 END RTL; --sinhw_altpriority_encoder_be8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altpriority_encoder_r08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END sinhw_altpriority_encoder_r08;

 ARCHITECTURE RTL OF sinhw_altpriority_encoder_r08 IS

	 SIGNAL  wire_altpriority_encoder5_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_w_lg_w_lg_zero12999w13000w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_w_lg_zero13001w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_w_lg_zero12999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_w_lg_w_lg_zero13001w13002w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_zero	:	STD_LOGIC;
	 COMPONENT  sinhw_altpriority_encoder_bv7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder6_w_lg_zero12999w & wire_altpriority_encoder6_w_lg_w_lg_zero13001w13002w);
	altpriority_encoder5 :  sinhw_altpriority_encoder_bv7
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder5_q
	  );
	loop44 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder6_w_lg_w_lg_zero12999w13000w(i) <= wire_altpriority_encoder6_w_lg_zero12999w(0) AND wire_altpriority_encoder6_q(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder6_w_lg_zero13001w(i) <= wire_altpriority_encoder6_zero AND wire_altpriority_encoder5_q(i);
	END GENERATE loop45;
	wire_altpriority_encoder6_w_lg_zero12999w(0) <= NOT wire_altpriority_encoder6_zero;
	loop46 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder6_w_lg_w_lg_zero13001w13002w(i) <= wire_altpriority_encoder6_w_lg_zero13001w(i) OR wire_altpriority_encoder6_w_lg_w_lg_zero12999w13000w(i);
	END GENERATE loop46;
	altpriority_encoder6 :  sinhw_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder6_q,
		zero => wire_altpriority_encoder6_zero
	  );

 END RTL; --sinhw_altpriority_encoder_r08


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altpriority_encoder_rf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END sinhw_altpriority_encoder_rf8;

 ARCHITECTURE RTL OF sinhw_altpriority_encoder_rf8 IS

	 SIGNAL  wire_altpriority_encoder15_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero13055w13056w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero13057w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero13055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero13057w13058w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_zero	:	STD_LOGIC;
	 COMPONENT  sinhw_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder16_w_lg_zero13055w & wire_altpriority_encoder16_w_lg_w_lg_zero13057w13058w);
	zero <= (wire_altpriority_encoder15_zero AND wire_altpriority_encoder16_zero);
	altpriority_encoder15 :  sinhw_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder15_q,
		zero => wire_altpriority_encoder15_zero
	  );
	loop47 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder16_w_lg_w_lg_zero13055w13056w(i) <= wire_altpriority_encoder16_w_lg_zero13055w(0) AND wire_altpriority_encoder16_q(i);
	END GENERATE loop47;
	loop48 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder16_w_lg_zero13057w(i) <= wire_altpriority_encoder16_zero AND wire_altpriority_encoder15_q(i);
	END GENERATE loop48;
	wire_altpriority_encoder16_w_lg_zero13055w(0) <= NOT wire_altpriority_encoder16_zero;
	loop49 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder16_w_lg_w_lg_zero13057w13058w(i) <= wire_altpriority_encoder16_w_lg_zero13057w(i) OR wire_altpriority_encoder16_w_lg_w_lg_zero13055w13056w(i);
	END GENERATE loop49;
	altpriority_encoder16 :  sinhw_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder16_q,
		zero => wire_altpriority_encoder16_zero
	  );

 END RTL; --sinhw_altpriority_encoder_rf8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altpriority_encoder_qb6 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END sinhw_altpriority_encoder_qb6;

 ARCHITECTURE RTL OF sinhw_altpriority_encoder_qb6 IS

	 SIGNAL  wire_altpriority_encoder3_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_w_lg_w_lg_zero12990w12991w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_w_lg_zero12992w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_w_lg_zero12990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_w_lg_w_lg_zero12992w12993w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_zero	:	STD_LOGIC;
	 COMPONENT  sinhw_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder4_w_lg_zero12990w & wire_altpriority_encoder4_w_lg_w_lg_zero12992w12993w);
	altpriority_encoder3 :  sinhw_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder3_q
	  );
	loop50 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder4_w_lg_w_lg_zero12990w12991w(i) <= wire_altpriority_encoder4_w_lg_zero12990w(0) AND wire_altpriority_encoder4_q(i);
	END GENERATE loop50;
	loop51 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder4_w_lg_zero12992w(i) <= wire_altpriority_encoder4_zero AND wire_altpriority_encoder3_q(i);
	END GENERATE loop51;
	wire_altpriority_encoder4_w_lg_zero12990w(0) <= NOT wire_altpriority_encoder4_zero;
	loop52 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder4_w_lg_w_lg_zero12992w12993w(i) <= wire_altpriority_encoder4_w_lg_zero12992w(i) OR wire_altpriority_encoder4_w_lg_w_lg_zero12990w12991w(i);
	END GENERATE loop52;
	altpriority_encoder4 :  sinhw_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder4_q,
		zero => wire_altpriority_encoder4_zero
	  );

 END RTL; --sinhw_altpriority_encoder_qb6

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 8 lpm_clshift 2 lpm_mult 1 lpm_mux 1 reg 780 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_range_b6c IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 circle	:	OUT  STD_LOGIC_VECTOR (35 DOWNTO 0);
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
		 negcircle	:	OUT  STD_LOGIC_VECTOR (35 DOWNTO 0)
	 ); 
 END sinhw_altfp_sincos_range_b6c;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_range_b6c IS

	 SIGNAL  wire_fp_range_table1_basefraction	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_fp_range_table1_incexponent	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_fp_range_table1_incmantissa	:	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  wire_clz23_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_clz23_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL	 basefractiondelff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 basefractionff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_0	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_1	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_2	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_3	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_4	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_5	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 circleff	:	STD_LOGIC_VECTOR(36 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponentff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 incexponentff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 incmantissaff	:	STD_LOGIC_VECTOR(55 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 leadff	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissadelff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissaff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissamultiplierff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 multipliernormff	:	STD_LOGIC_VECTOR(77 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 negbasefractiondelff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 negcircleff	:	STD_LOGIC_VECTOR(36 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 negrangeexponentff4	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 negrangeexponentff5	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_negrangeexponentff5_w_lg_w_lg_w_q_range11460w11464w11465w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_lg_w_q_range11460w11462w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_lg_w_q_range11460w11464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_q_range11461w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_q_range11460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rangeexponentff_0	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_1	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_2	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_3	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_4	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_5	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rangeexponentff_5_w_q_range11463w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 rotateff	:	STD_LOGIC_VECTOR(77 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rotateff_w_lg_w_q_range11477w11478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11481w11482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11484w11485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11487w11488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11490w11491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11493w11494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11496w11497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11499w11500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11502w11503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11505w11506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11508w11509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11511w11512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11514w11515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11517w11518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11520w11521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11523w11524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11526w11527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11529w11530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11532w11533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11535w11536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11538w11539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11541w11542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11544w11545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11547w11548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11550w11551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11553w11554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11556w11557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11559w11560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11562w11563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11565w11566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11568w11569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11571w11572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11574w11575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11577w11578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11580w11581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range11583w11584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range11583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 tableaddressff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_circle_add_dataa	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_circle_add_datab	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_circle_add_result	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_exponent_adjust_sub_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exponent_adjust_sub_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_negbasedractiondel_sub_dataa	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_negbasedractiondel_sub_result	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_negcircle_add_dataa	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_negcircle_add_datab	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_negcircle_add_result	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_negrangeexponent_sub4_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_negrangeexponent_sub4_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_negrangeexponent_sub5_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_negrangeexponent_sub5_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rangeexponent_sub1_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rangeexponent_sub1_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rangeexponent_sub5_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rangeexponent_sub5_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csftin_result	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_fp_lsft_rsft78_distance	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_lg_w_lg_w_lg_w_q_range11460w11464w11465w11466w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_fp_lsft_rsft78_result	:	STD_LOGIC_VECTOR (77 DOWNTO 0);
	 SIGNAL  wire_mult23x56_result	:	STD_LOGIC_VECTOR (78 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11069w11070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11117w11121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11117w11118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11122w11126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11122w11123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11127w11131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11127w11128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11132w11136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11132w11133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11137w11141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11137w11138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11142w11146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11142w11143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11147w11151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11147w11148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11152w11156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11152w11153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11157w11161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11157w11158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11162w11166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11162w11163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11071w11076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11071w11072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11167w11171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11167w11168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11172w11176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11172w11173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11177w11181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11177w11178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11182w11186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11182w11183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11187w11191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11187w11188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11192w11196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11192w11193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11197w11201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11197w11198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11202w11206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11202w11203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11207w11211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11207w11208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11212w11216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11212w11213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11077w11081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11077w11078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11217w11221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11217w11218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11222w11226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11222w11223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11227w11231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11227w11228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11232w11236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11232w11233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11237w11241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11237w11238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11242w11246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11242w11243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11247w11251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11247w11248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11252w11256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11252w11253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11257w11261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11257w11258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11262w11266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11262w11263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11082w11086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11082w11083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11267w11271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11267w11268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11272w11276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11272w11273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11277w11281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11277w11278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11282w11286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11282w11283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11287w11291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11287w11288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11292w11296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11292w11293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11297w11301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11297w11298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11302w11306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11302w11303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11307w11311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11307w11308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11312w11316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11312w11313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11087w11091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11087w11088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11317w11321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11317w11318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11322w11326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11322w11323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11327w11331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11327w11328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11332w11336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11332w11333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11337w11341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11337w11338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11342w11346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11342w11343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11347w11351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11347w11348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11352w11356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11352w11353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11357w11361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11357w11358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11362w11366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11362w11363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11092w11096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11092w11093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11367w11371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11367w11368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11372w11376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11372w11373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11377w11381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11377w11378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11382w11386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11382w11383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11387w11391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11387w11388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11392w11396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11392w11393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11397w11401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11397w11398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11402w11406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11402w11403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11407w11411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11407w11408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11412w11416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11412w11413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11097w11101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11097w11098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11417w11421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11417w11418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11422w11426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11422w11423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11427w11431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11427w11428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11432w11436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11432w11433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11437w11441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11437w11438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11442w11446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11442w11443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11447w11451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11447w11448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11452w11456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11452w11453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11102w11106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11102w11103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11107w11111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11107w11108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11112w11116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11112w11113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w11114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  basefractiondelnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  basefractionnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  circlenode_w :	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  const_23_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  incexponentnode_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  incmantissanode_w :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  leadnode_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  mantissaexponentnode_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  mantissamultipliernode_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  multipliernode_w :	STD_LOGIC_VECTOR (78 DOWNTO 0);
	 SIGNAL  multipliernormnode_w :	STD_LOGIC_VECTOR (77 DOWNTO 0);
	 SIGNAL  negbasefractiondelnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  negcirclenode_w :	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  negrotatenode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  rotatenode_w :	STD_LOGIC_VECTOR (77 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_data_range11039w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_data_range11040w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range11112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  sinhw_altfp_sincos_srrt_koa
	 PORT
	 ( 
		address	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		basefraction	:	OUT  STD_LOGIC_VECTOR(35 DOWNTO 0);
		incexponent	:	OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		incmantissa	:	OUT  STD_LOGIC_VECTOR(55 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altpriority_encoder_qb6
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_clshift
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_SHIFTTYPE	:	STRING := "LOGICAL";
		LPM_WIDTH	:	NATURAL;
		LPM_WIDTHDIST	:	NATURAL;
		lpm_type	:	STRING := "lpm_clshift"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		direction	:	IN STD_LOGIC := '0';
		distance	:	IN STD_LOGIC_VECTOR(LPM_WIDTHDIST-1 DOWNTO 0);
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		underflow	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11069w11070w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11069w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11117w11121w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11117w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11117w11118w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11117w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11122w11126w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11122w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11122w11123w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11122w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11127w11131w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11127w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11127w11128w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11127w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11132w11136w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11132w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11132w11133w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11132w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11137w11141w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11137w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11137w11138w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11137w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11142w11146w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11142w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11142w11143w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11142w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11147w11151w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11147w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11147w11148w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11147w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11152w11156w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11152w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11152w11153w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11152w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11157w11161w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11157w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11157w11158w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11157w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11162w11166w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11162w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11162w11163w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11162w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11071w11076w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11071w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11071w11072w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11071w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11167w11171w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11167w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11167w11168w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11167w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11172w11176w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11172w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11172w11173w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11172w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11177w11181w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11177w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11177w11178w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11177w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11182w11186w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11182w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11182w11183w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11182w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11187w11191w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11187w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11187w11188w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11187w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11192w11196w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11192w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11192w11193w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11192w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11197w11201w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11197w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11197w11198w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11197w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11202w11206w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11202w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11202w11203w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11202w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11207w11211w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11207w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11207w11208w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11207w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11212w11216w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11212w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11212w11213w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11212w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11077w11081w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11077w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11077w11078w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11077w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11217w11221w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11217w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11217w11218w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11217w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11222w11226w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11222w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11222w11223w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11222w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11227w11231w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11227w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11227w11228w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11227w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11232w11236w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11232w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11232w11233w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11232w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11237w11241w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11237w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11237w11238w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11237w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11242w11246w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11242w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11242w11243w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11242w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11247w11251w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11247w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11247w11248w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11247w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11252w11256w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11252w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11252w11253w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11252w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11257w11261w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11257w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11257w11258w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11257w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11262w11266w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11262w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11262w11263w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11262w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11082w11086w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11082w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11082w11083w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11082w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11267w11271w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11267w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11267w11268w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11267w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11272w11276w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11272w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11272w11273w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11272w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11277w11281w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11277w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11277w11278w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11277w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11282w11286w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11282w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11282w11283w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11282w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11287w11291w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11287w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11287w11288w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11287w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11292w11296w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11292w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11292w11293w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11292w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11297w11301w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11297w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11297w11298w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11297w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11302w11306w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11302w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11302w11303w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11302w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11307w11311w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11307w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11307w11308w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11307w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11312w11316w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11312w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11312w11313w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11312w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11087w11091w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11087w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11087w11088w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11087w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11317w11321w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11317w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11317w11318w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11317w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11322w11326w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11322w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11322w11323w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11322w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11327w11331w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11327w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11327w11328w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11327w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11332w11336w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11332w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11332w11333w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11332w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11337w11341w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11337w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11337w11338w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11337w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11342w11346w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11342w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11342w11343w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11342w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11347w11351w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11347w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11347w11348w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11347w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11352w11356w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11352w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11352w11353w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11352w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11357w11361w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11357w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11357w11358w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11357w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11362w11366w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11362w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11362w11363w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11362w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11092w11096w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11092w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11092w11093w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11092w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11367w11371w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11367w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11367w11368w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11367w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11372w11376w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11372w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11372w11373w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11372w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11377w11381w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11377w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11377w11378w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11377w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11382w11386w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11382w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11382w11383w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11382w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11387w11391w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11387w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11387w11388w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11387w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11392w11396w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11392w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11392w11393w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11392w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11397w11401w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11397w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11397w11398w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11397w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11402w11406w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11402w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11402w11403w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11402w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11407w11411w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11407w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11407w11408w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11407w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11412w11416w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11412w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11412w11413w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11412w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11097w11101w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11097w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11097w11098w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11097w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11417w11421w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11417w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11417w11418w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11417w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11422w11426w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11422w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11422w11423w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11422w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11427w11431w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11427w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11427w11428w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11427w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11432w11436w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11432w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11432w11433w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11432w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11437w11441w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11437w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11437w11438w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11437w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11442w11446w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11442w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11442w11443w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11442w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11447w11451w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11447w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11447w11448w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11447w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11452w11456w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11452w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11452w11453w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11452w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11457w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11048w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11102w11106w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11102w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11102w11103w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11102w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11107w11111w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11107w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11107w11108w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11107w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11112w11116w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11112w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11112w11113w(0) <= wire_crr_fp_range1_w_multipliernode_w_range11112w(0) AND wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w(0) <= NOT wire_crr_fp_range1_w_multipliernode_w_range11048w(0);
	wire_crr_fp_range1_w11119w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11117w11118w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11112w11116w(0);
	wire_crr_fp_range1_w11124w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11122w11123w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11117w11121w(0);
	wire_crr_fp_range1_w11129w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11127w11128w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11122w11126w(0);
	wire_crr_fp_range1_w11134w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11132w11133w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11127w11131w(0);
	wire_crr_fp_range1_w11139w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11137w11138w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11132w11136w(0);
	wire_crr_fp_range1_w11144w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11142w11143w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11137w11141w(0);
	wire_crr_fp_range1_w11149w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11147w11148w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11142w11146w(0);
	wire_crr_fp_range1_w11154w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11152w11153w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11147w11151w(0);
	wire_crr_fp_range1_w11159w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11157w11158w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11152w11156w(0);
	wire_crr_fp_range1_w11164w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11162w11163w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11157w11161w(0);
	wire_crr_fp_range1_w11073w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11071w11072w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11069w11070w(0);
	wire_crr_fp_range1_w11169w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11167w11168w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11162w11166w(0);
	wire_crr_fp_range1_w11174w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11172w11173w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11167w11171w(0);
	wire_crr_fp_range1_w11179w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11177w11178w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11172w11176w(0);
	wire_crr_fp_range1_w11184w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11182w11183w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11177w11181w(0);
	wire_crr_fp_range1_w11189w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11187w11188w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11182w11186w(0);
	wire_crr_fp_range1_w11194w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11192w11193w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11187w11191w(0);
	wire_crr_fp_range1_w11199w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11197w11198w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11192w11196w(0);
	wire_crr_fp_range1_w11204w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11202w11203w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11197w11201w(0);
	wire_crr_fp_range1_w11209w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11207w11208w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11202w11206w(0);
	wire_crr_fp_range1_w11214w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11212w11213w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11207w11211w(0);
	wire_crr_fp_range1_w11079w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11077w11078w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11071w11076w(0);
	wire_crr_fp_range1_w11219w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11217w11218w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11212w11216w(0);
	wire_crr_fp_range1_w11224w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11222w11223w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11217w11221w(0);
	wire_crr_fp_range1_w11229w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11227w11228w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11222w11226w(0);
	wire_crr_fp_range1_w11234w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11232w11233w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11227w11231w(0);
	wire_crr_fp_range1_w11239w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11237w11238w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11232w11236w(0);
	wire_crr_fp_range1_w11244w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11242w11243w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11237w11241w(0);
	wire_crr_fp_range1_w11249w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11247w11248w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11242w11246w(0);
	wire_crr_fp_range1_w11254w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11252w11253w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11247w11251w(0);
	wire_crr_fp_range1_w11259w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11257w11258w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11252w11256w(0);
	wire_crr_fp_range1_w11264w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11262w11263w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11257w11261w(0);
	wire_crr_fp_range1_w11084w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11082w11083w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11077w11081w(0);
	wire_crr_fp_range1_w11269w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11267w11268w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11262w11266w(0);
	wire_crr_fp_range1_w11274w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11272w11273w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11267w11271w(0);
	wire_crr_fp_range1_w11279w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11277w11278w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11272w11276w(0);
	wire_crr_fp_range1_w11284w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11282w11283w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11277w11281w(0);
	wire_crr_fp_range1_w11289w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11287w11288w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11282w11286w(0);
	wire_crr_fp_range1_w11294w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11292w11293w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11287w11291w(0);
	wire_crr_fp_range1_w11299w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11297w11298w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11292w11296w(0);
	wire_crr_fp_range1_w11304w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11302w11303w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11297w11301w(0);
	wire_crr_fp_range1_w11309w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11307w11308w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11302w11306w(0);
	wire_crr_fp_range1_w11314w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11312w11313w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11307w11311w(0);
	wire_crr_fp_range1_w11089w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11087w11088w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11082w11086w(0);
	wire_crr_fp_range1_w11319w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11317w11318w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11312w11316w(0);
	wire_crr_fp_range1_w11324w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11322w11323w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11317w11321w(0);
	wire_crr_fp_range1_w11329w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11327w11328w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11322w11326w(0);
	wire_crr_fp_range1_w11334w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11332w11333w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11327w11331w(0);
	wire_crr_fp_range1_w11339w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11337w11338w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11332w11336w(0);
	wire_crr_fp_range1_w11344w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11342w11343w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11337w11341w(0);
	wire_crr_fp_range1_w11349w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11347w11348w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11342w11346w(0);
	wire_crr_fp_range1_w11354w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11352w11353w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11347w11351w(0);
	wire_crr_fp_range1_w11359w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11357w11358w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11352w11356w(0);
	wire_crr_fp_range1_w11364w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11362w11363w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11357w11361w(0);
	wire_crr_fp_range1_w11094w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11092w11093w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11087w11091w(0);
	wire_crr_fp_range1_w11369w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11367w11368w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11362w11366w(0);
	wire_crr_fp_range1_w11374w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11372w11373w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11367w11371w(0);
	wire_crr_fp_range1_w11379w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11377w11378w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11372w11376w(0);
	wire_crr_fp_range1_w11384w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11382w11383w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11377w11381w(0);
	wire_crr_fp_range1_w11389w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11387w11388w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11382w11386w(0);
	wire_crr_fp_range1_w11394w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11392w11393w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11387w11391w(0);
	wire_crr_fp_range1_w11399w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11397w11398w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11392w11396w(0);
	wire_crr_fp_range1_w11404w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11402w11403w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11397w11401w(0);
	wire_crr_fp_range1_w11409w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11407w11408w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11402w11406w(0);
	wire_crr_fp_range1_w11414w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11412w11413w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11407w11411w(0);
	wire_crr_fp_range1_w11099w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11097w11098w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11092w11096w(0);
	wire_crr_fp_range1_w11419w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11417w11418w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11412w11416w(0);
	wire_crr_fp_range1_w11424w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11422w11423w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11417w11421w(0);
	wire_crr_fp_range1_w11429w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11427w11428w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11422w11426w(0);
	wire_crr_fp_range1_w11434w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11432w11433w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11427w11431w(0);
	wire_crr_fp_range1_w11439w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11437w11438w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11432w11436w(0);
	wire_crr_fp_range1_w11444w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11442w11443w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11437w11441w(0);
	wire_crr_fp_range1_w11449w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11447w11448w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11442w11446w(0);
	wire_crr_fp_range1_w11454w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11452w11453w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11447w11451w(0);
	wire_crr_fp_range1_w11458w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11457w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11452w11456w(0);
	wire_crr_fp_range1_w11104w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11102w11103w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11097w11101w(0);
	wire_crr_fp_range1_w11109w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11107w11108w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11102w11106w(0);
	wire_crr_fp_range1_w11114w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range11112w11113w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range11107w11111w(0);
	basefractiondelnode_w <= cbfd_5;
	basefractionnode_w <= wire_fp_range_table1_basefraction;
	circle <= circleff(35 DOWNTO 0);
	circlenode_w <= wire_circle_add_result;
	const_23_w <= "000010111";
	incexponentnode_w <= wire_fp_range_table1_incexponent;
	incmantissanode_w <= wire_fp_range_table1_incmantissa;
	leadnode_w <= (NOT wire_clz23_q);
	mantissaexponentnode_w <= wire_exponent_adjust_sub_result;
	mantissamultipliernode_w <= wire_csftin_result;
	multipliernode_w <= wire_mult23x56_result;
	multipliernormnode_w <= ( wire_crr_fp_range1_w11458w & wire_crr_fp_range1_w11454w & wire_crr_fp_range1_w11449w & wire_crr_fp_range1_w11444w & wire_crr_fp_range1_w11439w & wire_crr_fp_range1_w11434w & wire_crr_fp_range1_w11429w & wire_crr_fp_range1_w11424w & wire_crr_fp_range1_w11419w & wire_crr_fp_range1_w11414w & wire_crr_fp_range1_w11409w & wire_crr_fp_range1_w11404w & wire_crr_fp_range1_w11399w & wire_crr_fp_range1_w11394w & wire_crr_fp_range1_w11389w & wire_crr_fp_range1_w11384w & wire_crr_fp_range1_w11379w & wire_crr_fp_range1_w11374w & wire_crr_fp_range1_w11369w & wire_crr_fp_range1_w11364w & wire_crr_fp_range1_w11359w & wire_crr_fp_range1_w11354w & wire_crr_fp_range1_w11349w & wire_crr_fp_range1_w11344w & wire_crr_fp_range1_w11339w & wire_crr_fp_range1_w11334w & wire_crr_fp_range1_w11329w & wire_crr_fp_range1_w11324w & wire_crr_fp_range1_w11319w & wire_crr_fp_range1_w11314w & wire_crr_fp_range1_w11309w & wire_crr_fp_range1_w11304w & wire_crr_fp_range1_w11299w & wire_crr_fp_range1_w11294w & wire_crr_fp_range1_w11289w & wire_crr_fp_range1_w11284w & wire_crr_fp_range1_w11279w & wire_crr_fp_range1_w11274w & wire_crr_fp_range1_w11269w & wire_crr_fp_range1_w11264w & wire_crr_fp_range1_w11259w & wire_crr_fp_range1_w11254w & wire_crr_fp_range1_w11249w & wire_crr_fp_range1_w11244w & wire_crr_fp_range1_w11239w & wire_crr_fp_range1_w11234w & wire_crr_fp_range1_w11229w & wire_crr_fp_range1_w11224w & wire_crr_fp_range1_w11219w & wire_crr_fp_range1_w11214w & wire_crr_fp_range1_w11209w & wire_crr_fp_range1_w11204w & wire_crr_fp_range1_w11199w & wire_crr_fp_range1_w11194w & wire_crr_fp_range1_w11189w & wire_crr_fp_range1_w11184w & wire_crr_fp_range1_w11179w & wire_crr_fp_range1_w11174w & wire_crr_fp_range1_w11169w & wire_crr_fp_range1_w11164w & wire_crr_fp_range1_w11159w & wire_crr_fp_range1_w11154w & wire_crr_fp_range1_w11149w & wire_crr_fp_range1_w11144w & wire_crr_fp_range1_w11139w & wire_crr_fp_range1_w11134w & wire_crr_fp_range1_w11129w & wire_crr_fp_range1_w11124w & wire_crr_fp_range1_w11119w & wire_crr_fp_range1_w11114w
 & wire_crr_fp_range1_w11109w & wire_crr_fp_range1_w11104w & wire_crr_fp_range1_w11099w & wire_crr_fp_range1_w11094w & wire_crr_fp_range1_w11089w & wire_crr_fp_range1_w11084w & wire_crr_fp_range1_w11079w & wire_crr_fp_range1_w11073w);
	negbasefractiondelnode_w <= wire_negbasedractiondel_sub_result;
	negcircle <= negcircleff(35 DOWNTO 0);
	negcirclenode_w <= wire_negcircle_add_result;
	negrotatenode_w <= ( wire_rotateff_w_lg_w_q_range11583w11584w & wire_rotateff_w_lg_w_q_range11580w11581w & wire_rotateff_w_lg_w_q_range11577w11578w & wire_rotateff_w_lg_w_q_range11574w11575w & wire_rotateff_w_lg_w_q_range11571w11572w & wire_rotateff_w_lg_w_q_range11568w11569w & wire_rotateff_w_lg_w_q_range11565w11566w & wire_rotateff_w_lg_w_q_range11562w11563w & wire_rotateff_w_lg_w_q_range11559w11560w & wire_rotateff_w_lg_w_q_range11556w11557w & wire_rotateff_w_lg_w_q_range11553w11554w & wire_rotateff_w_lg_w_q_range11550w11551w & wire_rotateff_w_lg_w_q_range11547w11548w & wire_rotateff_w_lg_w_q_range11544w11545w & wire_rotateff_w_lg_w_q_range11541w11542w & wire_rotateff_w_lg_w_q_range11538w11539w & wire_rotateff_w_lg_w_q_range11535w11536w & wire_rotateff_w_lg_w_q_range11532w11533w & wire_rotateff_w_lg_w_q_range11529w11530w & wire_rotateff_w_lg_w_q_range11526w11527w & wire_rotateff_w_lg_w_q_range11523w11524w & wire_rotateff_w_lg_w_q_range11520w11521w & wire_rotateff_w_lg_w_q_range11517w11518w & wire_rotateff_w_lg_w_q_range11514w11515w & wire_rotateff_w_lg_w_q_range11511w11512w & wire_rotateff_w_lg_w_q_range11508w11509w & wire_rotateff_w_lg_w_q_range11505w11506w & wire_rotateff_w_lg_w_q_range11502w11503w & wire_rotateff_w_lg_w_q_range11499w11500w & wire_rotateff_w_lg_w_q_range11496w11497w & wire_rotateff_w_lg_w_q_range11493w11494w & wire_rotateff_w_lg_w_q_range11490w11491w & wire_rotateff_w_lg_w_q_range11487w11488w & wire_rotateff_w_lg_w_q_range11484w11485w & wire_rotateff_w_lg_w_q_range11481w11482w & wire_rotateff_w_lg_w_q_range11477w11478w);
	rotatenode_w <= wire_fp_lsft_rsft78_result;
	wire_crr_fp_range1_w_data_range11039w <= data(22 DOWNTO 0);
	wire_crr_fp_range1_w_data_range11040w <= data(30 DOWNTO 23);
	wire_crr_fp_range1_w_multipliernode_w_range11069w(0) <= multipliernode_w(0);
	wire_crr_fp_range1_w_multipliernode_w_range11117w(0) <= multipliernode_w(10);
	wire_crr_fp_range1_w_multipliernode_w_range11122w(0) <= multipliernode_w(11);
	wire_crr_fp_range1_w_multipliernode_w_range11127w(0) <= multipliernode_w(12);
	wire_crr_fp_range1_w_multipliernode_w_range11132w(0) <= multipliernode_w(13);
	wire_crr_fp_range1_w_multipliernode_w_range11137w(0) <= multipliernode_w(14);
	wire_crr_fp_range1_w_multipliernode_w_range11142w(0) <= multipliernode_w(15);
	wire_crr_fp_range1_w_multipliernode_w_range11147w(0) <= multipliernode_w(16);
	wire_crr_fp_range1_w_multipliernode_w_range11152w(0) <= multipliernode_w(17);
	wire_crr_fp_range1_w_multipliernode_w_range11157w(0) <= multipliernode_w(18);
	wire_crr_fp_range1_w_multipliernode_w_range11162w(0) <= multipliernode_w(19);
	wire_crr_fp_range1_w_multipliernode_w_range11071w(0) <= multipliernode_w(1);
	wire_crr_fp_range1_w_multipliernode_w_range11167w(0) <= multipliernode_w(20);
	wire_crr_fp_range1_w_multipliernode_w_range11172w(0) <= multipliernode_w(21);
	wire_crr_fp_range1_w_multipliernode_w_range11177w(0) <= multipliernode_w(22);
	wire_crr_fp_range1_w_multipliernode_w_range11182w(0) <= multipliernode_w(23);
	wire_crr_fp_range1_w_multipliernode_w_range11187w(0) <= multipliernode_w(24);
	wire_crr_fp_range1_w_multipliernode_w_range11192w(0) <= multipliernode_w(25);
	wire_crr_fp_range1_w_multipliernode_w_range11197w(0) <= multipliernode_w(26);
	wire_crr_fp_range1_w_multipliernode_w_range11202w(0) <= multipliernode_w(27);
	wire_crr_fp_range1_w_multipliernode_w_range11207w(0) <= multipliernode_w(28);
	wire_crr_fp_range1_w_multipliernode_w_range11212w(0) <= multipliernode_w(29);
	wire_crr_fp_range1_w_multipliernode_w_range11077w(0) <= multipliernode_w(2);
	wire_crr_fp_range1_w_multipliernode_w_range11217w(0) <= multipliernode_w(30);
	wire_crr_fp_range1_w_multipliernode_w_range11222w(0) <= multipliernode_w(31);
	wire_crr_fp_range1_w_multipliernode_w_range11227w(0) <= multipliernode_w(32);
	wire_crr_fp_range1_w_multipliernode_w_range11232w(0) <= multipliernode_w(33);
	wire_crr_fp_range1_w_multipliernode_w_range11237w(0) <= multipliernode_w(34);
	wire_crr_fp_range1_w_multipliernode_w_range11242w(0) <= multipliernode_w(35);
	wire_crr_fp_range1_w_multipliernode_w_range11247w(0) <= multipliernode_w(36);
	wire_crr_fp_range1_w_multipliernode_w_range11252w(0) <= multipliernode_w(37);
	wire_crr_fp_range1_w_multipliernode_w_range11257w(0) <= multipliernode_w(38);
	wire_crr_fp_range1_w_multipliernode_w_range11262w(0) <= multipliernode_w(39);
	wire_crr_fp_range1_w_multipliernode_w_range11082w(0) <= multipliernode_w(3);
	wire_crr_fp_range1_w_multipliernode_w_range11267w(0) <= multipliernode_w(40);
	wire_crr_fp_range1_w_multipliernode_w_range11272w(0) <= multipliernode_w(41);
	wire_crr_fp_range1_w_multipliernode_w_range11277w(0) <= multipliernode_w(42);
	wire_crr_fp_range1_w_multipliernode_w_range11282w(0) <= multipliernode_w(43);
	wire_crr_fp_range1_w_multipliernode_w_range11287w(0) <= multipliernode_w(44);
	wire_crr_fp_range1_w_multipliernode_w_range11292w(0) <= multipliernode_w(45);
	wire_crr_fp_range1_w_multipliernode_w_range11297w(0) <= multipliernode_w(46);
	wire_crr_fp_range1_w_multipliernode_w_range11302w(0) <= multipliernode_w(47);
	wire_crr_fp_range1_w_multipliernode_w_range11307w(0) <= multipliernode_w(48);
	wire_crr_fp_range1_w_multipliernode_w_range11312w(0) <= multipliernode_w(49);
	wire_crr_fp_range1_w_multipliernode_w_range11087w(0) <= multipliernode_w(4);
	wire_crr_fp_range1_w_multipliernode_w_range11317w(0) <= multipliernode_w(50);
	wire_crr_fp_range1_w_multipliernode_w_range11322w(0) <= multipliernode_w(51);
	wire_crr_fp_range1_w_multipliernode_w_range11327w(0) <= multipliernode_w(52);
	wire_crr_fp_range1_w_multipliernode_w_range11332w(0) <= multipliernode_w(53);
	wire_crr_fp_range1_w_multipliernode_w_range11337w(0) <= multipliernode_w(54);
	wire_crr_fp_range1_w_multipliernode_w_range11342w(0) <= multipliernode_w(55);
	wire_crr_fp_range1_w_multipliernode_w_range11347w(0) <= multipliernode_w(56);
	wire_crr_fp_range1_w_multipliernode_w_range11352w(0) <= multipliernode_w(57);
	wire_crr_fp_range1_w_multipliernode_w_range11357w(0) <= multipliernode_w(58);
	wire_crr_fp_range1_w_multipliernode_w_range11362w(0) <= multipliernode_w(59);
	wire_crr_fp_range1_w_multipliernode_w_range11092w(0) <= multipliernode_w(5);
	wire_crr_fp_range1_w_multipliernode_w_range11367w(0) <= multipliernode_w(60);
	wire_crr_fp_range1_w_multipliernode_w_range11372w(0) <= multipliernode_w(61);
	wire_crr_fp_range1_w_multipliernode_w_range11377w(0) <= multipliernode_w(62);
	wire_crr_fp_range1_w_multipliernode_w_range11382w(0) <= multipliernode_w(63);
	wire_crr_fp_range1_w_multipliernode_w_range11387w(0) <= multipliernode_w(64);
	wire_crr_fp_range1_w_multipliernode_w_range11392w(0) <= multipliernode_w(65);
	wire_crr_fp_range1_w_multipliernode_w_range11397w(0) <= multipliernode_w(66);
	wire_crr_fp_range1_w_multipliernode_w_range11402w(0) <= multipliernode_w(67);
	wire_crr_fp_range1_w_multipliernode_w_range11407w(0) <= multipliernode_w(68);
	wire_crr_fp_range1_w_multipliernode_w_range11412w(0) <= multipliernode_w(69);
	wire_crr_fp_range1_w_multipliernode_w_range11097w(0) <= multipliernode_w(6);
	wire_crr_fp_range1_w_multipliernode_w_range11417w(0) <= multipliernode_w(70);
	wire_crr_fp_range1_w_multipliernode_w_range11422w(0) <= multipliernode_w(71);
	wire_crr_fp_range1_w_multipliernode_w_range11427w(0) <= multipliernode_w(72);
	wire_crr_fp_range1_w_multipliernode_w_range11432w(0) <= multipliernode_w(73);
	wire_crr_fp_range1_w_multipliernode_w_range11437w(0) <= multipliernode_w(74);
	wire_crr_fp_range1_w_multipliernode_w_range11442w(0) <= multipliernode_w(75);
	wire_crr_fp_range1_w_multipliernode_w_range11447w(0) <= multipliernode_w(76);
	wire_crr_fp_range1_w_multipliernode_w_range11452w(0) <= multipliernode_w(77);
	wire_crr_fp_range1_w_multipliernode_w_range11048w(0) <= multipliernode_w(78);
	wire_crr_fp_range1_w_multipliernode_w_range11102w(0) <= multipliernode_w(7);
	wire_crr_fp_range1_w_multipliernode_w_range11107w(0) <= multipliernode_w(8);
	wire_crr_fp_range1_w_multipliernode_w_range11112w(0) <= multipliernode_w(9);
	fp_range_table1 :  sinhw_altfp_sincos_srrt_koa
	  PORT MAP ( 
		address => tableaddressff,
		basefraction => wire_fp_range_table1_basefraction,
		incexponent => wire_fp_range_table1_incexponent,
		incmantissa => wire_fp_range_table1_incmantissa
	  );
	wire_clz23_data <= ( mantissaff & "111111111");
	clz23 :  sinhw_altpriority_encoder_qb6
	  PORT MAP ( 
		data => wire_clz23_data,
		q => wire_clz23_q
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN basefractiondelff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN basefractiondelff <= basefractiondelnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN basefractionff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN basefractionff <= basefractionnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_0 <= basefractionff;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_1 <= cbfd_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_2 <= cbfd_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_3 <= cbfd_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_4 <= cbfd_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_5 <= cbfd_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN circleff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN circleff <= circlenode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponentff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN exponentff <= wire_crr_fp_range1_w_data_range11040w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN incexponentff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN incexponentff <= incexponentnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN incmantissaff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN incmantissaff <= incmantissanode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN leadff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN leadff <= leadnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissadelff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN mantissadelff <= mantissaff;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissaff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN mantissaff <= wire_crr_fp_range1_w_data_range11039w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissamultiplierff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN mantissamultiplierff <= mantissamultipliernode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN multipliernormff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN multipliernormff <= multipliernormnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN negbasefractiondelff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN negbasefractiondelff <= negbasefractiondelnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN negcircleff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN negcircleff <= negcirclenode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN negrangeexponentff4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN negrangeexponentff4 <= wire_negrangeexponent_sub4_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN negrangeexponentff5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN negrangeexponentff5 <= wire_negrangeexponent_sub5_result;
			END IF;
		END IF;
	END PROCESS;
	loop53 : FOR i IN 0 TO 6 GENERATE 
		wire_negrangeexponentff5_w_lg_w_lg_w_q_range11460w11464w11465w(i) <= wire_negrangeexponentff5_w_lg_w_q_range11460w11464w(0) AND wire_rangeexponentff_5_w_q_range11463w(i);
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 6 GENERATE 
		wire_negrangeexponentff5_w_lg_w_q_range11460w11462w(i) <= wire_negrangeexponentff5_w_q_range11460w(0) AND wire_negrangeexponentff5_w_q_range11461w(i);
	END GENERATE loop54;
	wire_negrangeexponentff5_w_lg_w_q_range11460w11464w(0) <= NOT wire_negrangeexponentff5_w_q_range11460w(0);
	wire_negrangeexponentff5_w_q_range11461w <= negrangeexponentff5(6 DOWNTO 0);
	wire_negrangeexponentff5_w_q_range11460w(0) <= negrangeexponentff5(8);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_0 <= mantissaexponentnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_1 <= wire_rangeexponent_sub1_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_2 <= rangeexponentff_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_3 <= rangeexponentff_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_4 <= rangeexponentff_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_5 <= wire_rangeexponent_sub5_result;
			END IF;
		END IF;
	END PROCESS;
	wire_rangeexponentff_5_w_q_range11463w <= rangeexponentff_5(6 DOWNTO 0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rotateff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rotateff <= rotatenode_w;
			END IF;
		END IF;
	END PROCESS;
	wire_rotateff_w_lg_w_q_range11477w11478w(0) <= NOT wire_rotateff_w_q_range11477w(0);
	wire_rotateff_w_lg_w_q_range11481w11482w(0) <= NOT wire_rotateff_w_q_range11481w(0);
	wire_rotateff_w_lg_w_q_range11484w11485w(0) <= NOT wire_rotateff_w_q_range11484w(0);
	wire_rotateff_w_lg_w_q_range11487w11488w(0) <= NOT wire_rotateff_w_q_range11487w(0);
	wire_rotateff_w_lg_w_q_range11490w11491w(0) <= NOT wire_rotateff_w_q_range11490w(0);
	wire_rotateff_w_lg_w_q_range11493w11494w(0) <= NOT wire_rotateff_w_q_range11493w(0);
	wire_rotateff_w_lg_w_q_range11496w11497w(0) <= NOT wire_rotateff_w_q_range11496w(0);
	wire_rotateff_w_lg_w_q_range11499w11500w(0) <= NOT wire_rotateff_w_q_range11499w(0);
	wire_rotateff_w_lg_w_q_range11502w11503w(0) <= NOT wire_rotateff_w_q_range11502w(0);
	wire_rotateff_w_lg_w_q_range11505w11506w(0) <= NOT wire_rotateff_w_q_range11505w(0);
	wire_rotateff_w_lg_w_q_range11508w11509w(0) <= NOT wire_rotateff_w_q_range11508w(0);
	wire_rotateff_w_lg_w_q_range11511w11512w(0) <= NOT wire_rotateff_w_q_range11511w(0);
	wire_rotateff_w_lg_w_q_range11514w11515w(0) <= NOT wire_rotateff_w_q_range11514w(0);
	wire_rotateff_w_lg_w_q_range11517w11518w(0) <= NOT wire_rotateff_w_q_range11517w(0);
	wire_rotateff_w_lg_w_q_range11520w11521w(0) <= NOT wire_rotateff_w_q_range11520w(0);
	wire_rotateff_w_lg_w_q_range11523w11524w(0) <= NOT wire_rotateff_w_q_range11523w(0);
	wire_rotateff_w_lg_w_q_range11526w11527w(0) <= NOT wire_rotateff_w_q_range11526w(0);
	wire_rotateff_w_lg_w_q_range11529w11530w(0) <= NOT wire_rotateff_w_q_range11529w(0);
	wire_rotateff_w_lg_w_q_range11532w11533w(0) <= NOT wire_rotateff_w_q_range11532w(0);
	wire_rotateff_w_lg_w_q_range11535w11536w(0) <= NOT wire_rotateff_w_q_range11535w(0);
	wire_rotateff_w_lg_w_q_range11538w11539w(0) <= NOT wire_rotateff_w_q_range11538w(0);
	wire_rotateff_w_lg_w_q_range11541w11542w(0) <= NOT wire_rotateff_w_q_range11541w(0);
	wire_rotateff_w_lg_w_q_range11544w11545w(0) <= NOT wire_rotateff_w_q_range11544w(0);
	wire_rotateff_w_lg_w_q_range11547w11548w(0) <= NOT wire_rotateff_w_q_range11547w(0);
	wire_rotateff_w_lg_w_q_range11550w11551w(0) <= NOT wire_rotateff_w_q_range11550w(0);
	wire_rotateff_w_lg_w_q_range11553w11554w(0) <= NOT wire_rotateff_w_q_range11553w(0);
	wire_rotateff_w_lg_w_q_range11556w11557w(0) <= NOT wire_rotateff_w_q_range11556w(0);
	wire_rotateff_w_lg_w_q_range11559w11560w(0) <= NOT wire_rotateff_w_q_range11559w(0);
	wire_rotateff_w_lg_w_q_range11562w11563w(0) <= NOT wire_rotateff_w_q_range11562w(0);
	wire_rotateff_w_lg_w_q_range11565w11566w(0) <= NOT wire_rotateff_w_q_range11565w(0);
	wire_rotateff_w_lg_w_q_range11568w11569w(0) <= NOT wire_rotateff_w_q_range11568w(0);
	wire_rotateff_w_lg_w_q_range11571w11572w(0) <= NOT wire_rotateff_w_q_range11571w(0);
	wire_rotateff_w_lg_w_q_range11574w11575w(0) <= NOT wire_rotateff_w_q_range11574w(0);
	wire_rotateff_w_lg_w_q_range11577w11578w(0) <= NOT wire_rotateff_w_q_range11577w(0);
	wire_rotateff_w_lg_w_q_range11580w11581w(0) <= NOT wire_rotateff_w_q_range11580w(0);
	wire_rotateff_w_lg_w_q_range11583w11584w(0) <= NOT wire_rotateff_w_q_range11583w(0);
	wire_rotateff_w_q_range11477w(0) <= rotateff(42);
	wire_rotateff_w_q_range11481w(0) <= rotateff(43);
	wire_rotateff_w_q_range11484w(0) <= rotateff(44);
	wire_rotateff_w_q_range11487w(0) <= rotateff(45);
	wire_rotateff_w_q_range11490w(0) <= rotateff(46);
	wire_rotateff_w_q_range11493w(0) <= rotateff(47);
	wire_rotateff_w_q_range11496w(0) <= rotateff(48);
	wire_rotateff_w_q_range11499w(0) <= rotateff(49);
	wire_rotateff_w_q_range11502w(0) <= rotateff(50);
	wire_rotateff_w_q_range11505w(0) <= rotateff(51);
	wire_rotateff_w_q_range11508w(0) <= rotateff(52);
	wire_rotateff_w_q_range11511w(0) <= rotateff(53);
	wire_rotateff_w_q_range11514w(0) <= rotateff(54);
	wire_rotateff_w_q_range11517w(0) <= rotateff(55);
	wire_rotateff_w_q_range11520w(0) <= rotateff(56);
	wire_rotateff_w_q_range11523w(0) <= rotateff(57);
	wire_rotateff_w_q_range11526w(0) <= rotateff(58);
	wire_rotateff_w_q_range11529w(0) <= rotateff(59);
	wire_rotateff_w_q_range11532w(0) <= rotateff(60);
	wire_rotateff_w_q_range11535w(0) <= rotateff(61);
	wire_rotateff_w_q_range11538w(0) <= rotateff(62);
	wire_rotateff_w_q_range11541w(0) <= rotateff(63);
	wire_rotateff_w_q_range11544w(0) <= rotateff(64);
	wire_rotateff_w_q_range11547w(0) <= rotateff(65);
	wire_rotateff_w_q_range11550w(0) <= rotateff(66);
	wire_rotateff_w_q_range11553w(0) <= rotateff(67);
	wire_rotateff_w_q_range11556w(0) <= rotateff(68);
	wire_rotateff_w_q_range11559w(0) <= rotateff(69);
	wire_rotateff_w_q_range11562w(0) <= rotateff(70);
	wire_rotateff_w_q_range11565w(0) <= rotateff(71);
	wire_rotateff_w_q_range11568w(0) <= rotateff(72);
	wire_rotateff_w_q_range11571w(0) <= rotateff(73);
	wire_rotateff_w_q_range11574w(0) <= rotateff(74);
	wire_rotateff_w_q_range11577w(0) <= rotateff(75);
	wire_rotateff_w_q_range11580w(0) <= rotateff(76);
	wire_rotateff_w_q_range11583w(0) <= rotateff(77);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tableaddressff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN tableaddressff <= exponentff;
			END IF;
		END IF;
	END PROCESS;
	wire_circle_add_dataa <= ( "0" & basefractiondelff);
	wire_circle_add_datab <= ( "0" & rotateff(77 DOWNTO 42));
	circle_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 37
	  )
	  PORT MAP ( 
		dataa => wire_circle_add_dataa,
		datab => wire_circle_add_datab,
		result => wire_circle_add_result
	  );
	wire_exponent_adjust_sub_datab <= ( "0000" & leadff);
	exponent_adjust_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => const_23_w,
		datab => wire_exponent_adjust_sub_datab,
		result => wire_exponent_adjust_sub_result
	  );
	wire_negbasedractiondel_sub_dataa <= (OTHERS => '0');
	negbasedractiondel_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 36
	  )
	  PORT MAP ( 
		dataa => wire_negbasedractiondel_sub_dataa,
		datab => basefractiondelnode_w(35 DOWNTO 0),
		result => wire_negbasedractiondel_sub_result
	  );
	wire_negcircle_add_dataa <= ( "1" & negbasefractiondelff);
	wire_negcircle_add_datab <= ( "1" & negrotatenode_w);
	negcircle_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 37
	  )
	  PORT MAP ( 
		cin => wire_vcc,
		dataa => wire_negcircle_add_dataa,
		datab => wire_negcircle_add_datab,
		result => wire_negcircle_add_result
	  );
	wire_negrangeexponent_sub4_dataa <= ( "1" & "00000000");
	negrangeexponent_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => wire_negrangeexponent_sub4_dataa,
		datab => rangeexponentff_3,
		result => wire_negrangeexponent_sub4_result
	  );
	wire_negrangeexponent_sub5_datab <= ( "00000000" & wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w);
	negrangeexponent_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => negrangeexponentff4,
		datab => wire_negrangeexponent_sub5_datab,
		result => wire_negrangeexponent_sub5_result
	  );
	wire_rangeexponent_sub1_datab <= ( "0" & incexponentff);
	rangeexponent_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => rangeexponentff_0,
		datab => wire_rangeexponent_sub1_datab,
		result => wire_rangeexponent_sub1_result
	  );
	wire_rangeexponent_sub5_datab <= ( "00000000" & wire_crr_fp_range1_w_lg_w_multipliernode_w_range11048w11049w);
	rangeexponent_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => rangeexponentff_4,
		datab => wire_rangeexponent_sub5_datab,
		result => wire_rangeexponent_sub5_result
	  );
	csftin :  lpm_clshift
	  GENERIC MAP (
		LPM_WIDTH => 23,
		LPM_WIDTHDIST => 5
	  )
	  PORT MAP ( 
		data => mantissadelff,
		direction => wire_gnd,
		distance => leadff,
		result => wire_csftin_result
	  );
	wire_fp_lsft_rsft78_distance <= wire_negrangeexponentff5_w_lg_w_lg_w_lg_w_q_range11460w11464w11465w11466w;
	loop55 : FOR i IN 0 TO 6 GENERATE 
		wire_negrangeexponentff5_w_lg_w_lg_w_lg_w_q_range11460w11464w11465w11466w(i) <= wire_negrangeexponentff5_w_lg_w_lg_w_q_range11460w11464w11465w(i) OR wire_negrangeexponentff5_w_lg_w_q_range11460w11462w(i);
	END GENERATE loop55;
	fp_lsft_rsft78 :  lpm_clshift
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_WIDTH => 78,
		LPM_WIDTHDIST => 7
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		data => multipliernormff,
		direction => negrangeexponentff5(8),
		distance => wire_fp_lsft_rsft78_distance,
		result => wire_fp_lsft_rsft78_result
	  );
	mult23x56 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 4,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 23,
		LPM_WIDTHB => 56,
		LPM_WIDTHP => 79
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => mantissamultiplierff,
		datab => incmantissaff,
		result => wire_mult23x56_result
	  );

 END RTL; --sinhw_altfp_sincos_range_b6c


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" WIDTH=64 WIDTHAD=6 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altpriority_encoder_q08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END sinhw_altpriority_encoder_q08;

 ARCHITECTURE RTL OF sinhw_altpriority_encoder_q08 IS

	 SIGNAL  wire_altpriority_encoder19_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero13074w13075w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero13076w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero13074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero13076w13077w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_zero	:	STD_LOGIC;
	 COMPONENT  sinhw_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder20_w_lg_zero13074w & wire_altpriority_encoder20_w_lg_w_lg_zero13076w13077w);
	altpriority_encoder19 :  sinhw_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder19_q
	  );
	loop56 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero13074w13075w(i) <= wire_altpriority_encoder20_w_lg_zero13074w(0) AND wire_altpriority_encoder20_q(i);
	END GENERATE loop56;
	loop57 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder20_w_lg_zero13076w(i) <= wire_altpriority_encoder20_zero AND wire_altpriority_encoder19_q(i);
	END GENERATE loop57;
	wire_altpriority_encoder20_w_lg_zero13074w(0) <= NOT wire_altpriority_encoder20_zero;
	loop58 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero13076w13077w(i) <= wire_altpriority_encoder20_w_lg_zero13076w(i) OR wire_altpriority_encoder20_w_lg_w_lg_zero13074w13075w(i);
	END GENERATE loop58;
	altpriority_encoder20 :  sinhw_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder20_q,
		zero => wire_altpriority_encoder20_zero
	  );

 END RTL; --sinhw_altpriority_encoder_q08


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=32 WIDTHAD=5 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altpriority_encoder_qf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END sinhw_altpriority_encoder_qf8;

 ARCHITECTURE RTL OF sinhw_altpriority_encoder_qf8 IS

	 SIGNAL  wire_altpriority_encoder21_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero13083w13084w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero13085w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero13083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero13085w13086w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_zero	:	STD_LOGIC;
	 COMPONENT  sinhw_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder22_w_lg_zero13083w & wire_altpriority_encoder22_w_lg_w_lg_zero13085w13086w);
	zero <= (wire_altpriority_encoder21_zero AND wire_altpriority_encoder22_zero);
	altpriority_encoder21 :  sinhw_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder21_q,
		zero => wire_altpriority_encoder21_zero
	  );
	loop59 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder22_w_lg_w_lg_zero13083w13084w(i) <= wire_altpriority_encoder22_w_lg_zero13083w(0) AND wire_altpriority_encoder22_q(i);
	END GENERATE loop59;
	loop60 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder22_w_lg_zero13085w(i) <= wire_altpriority_encoder22_zero AND wire_altpriority_encoder21_q(i);
	END GENERATE loop60;
	wire_altpriority_encoder22_w_lg_zero13083w(0) <= NOT wire_altpriority_encoder22_zero;
	loop61 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder22_w_lg_w_lg_zero13085w13086w(i) <= wire_altpriority_encoder22_w_lg_zero13085w(i) OR wire_altpriority_encoder22_w_lg_w_lg_zero13083w13084w(i);
	END GENERATE loop61;
	altpriority_encoder22 :  sinhw_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder22_q,
		zero => wire_altpriority_encoder22_zero
	  );

 END RTL; --sinhw_altpriority_encoder_qf8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altpriority_encoder_0c6 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0)
	 ); 
 END sinhw_altpriority_encoder_0c6;

 ARCHITECTURE RTL OF sinhw_altpriority_encoder_0c6 IS

	 SIGNAL  wire_altpriority_encoder17_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero13065w13066w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero13067w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero13065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero13067w13068w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_zero	:	STD_LOGIC;
	 COMPONENT  sinhw_altpriority_encoder_q08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altpriority_encoder_qf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder18_w_lg_zero13065w & wire_altpriority_encoder18_w_lg_w_lg_zero13067w13068w);
	altpriority_encoder17 :  sinhw_altpriority_encoder_q08
	  PORT MAP ( 
		data => data(31 DOWNTO 0),
		q => wire_altpriority_encoder17_q
	  );
	loop62 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder18_w_lg_w_lg_zero13065w13066w(i) <= wire_altpriority_encoder18_w_lg_zero13065w(0) AND wire_altpriority_encoder18_q(i);
	END GENERATE loop62;
	loop63 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder18_w_lg_zero13067w(i) <= wire_altpriority_encoder18_zero AND wire_altpriority_encoder17_q(i);
	END GENERATE loop63;
	wire_altpriority_encoder18_w_lg_zero13065w(0) <= NOT wire_altpriority_encoder18_zero;
	loop64 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder18_w_lg_w_lg_zero13067w13068w(i) <= wire_altpriority_encoder18_w_lg_zero13067w(i) OR wire_altpriority_encoder18_w_lg_w_lg_zero13065w13066w(i);
	END GENERATE loop64;
	altpriority_encoder18 :  sinhw_altpriority_encoder_qf8
	  PORT MAP ( 
		data => data(63 DOWNTO 32),
		q => wire_altpriority_encoder18_q,
		zero => wire_altpriority_encoder18_zero
	  );

 END RTL; --sinhw_altpriority_encoder_0c6

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 52 lpm_clshift 3 lpm_mult 3 lpm_mux 2 reg 3720 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  sinhw_altfp_sincos_47e IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END sinhw_altfp_sincos_47e;

 ARCHITECTURE RTL OF sinhw_altfp_sincos_47e IS

	 SIGNAL  wire_ccc_cordic_m_sincos	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_circle	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_negcircle	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_clz_data	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_clz_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL	 countff	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponentinff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponentnormff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exponentnormff_w_lg_q398w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exponentnormff_w_lg_w_lg_q398w399w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	 exponentoutff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 fixed_sincosff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_0	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_1	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_10	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_11	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_12	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_13	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_14	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_15	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_16	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_17	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_18	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_19	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_2	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_20	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_21	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_22	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_23	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_24	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_25	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_26	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_27	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_28	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_29	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_3	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_30	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_31	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_32	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_33	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_34	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_4	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_5	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_6	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_7	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_8	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 input_delay_ff_9	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissanormff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_mantissanormff_w_lg_q394w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_mantissanormff_w_lg_w_lg_q394w395w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL	 mantissaoutff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 quadrant_sumff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 select_sincosff	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 selectoutputff	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_selectoutputff_w_lg_w_q_range390w393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_selectoutputff_w_q_range390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 signcalcff	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_signcalcff_w_lg_w_q_range402w403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_signcalcff_w_q_range402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 signinff	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_signinff_w_q_range56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 signoutff	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exponentcheck_sub_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exponentcheck_sub_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exponentcheck_sub_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exponentnorm_add_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exponentnorm_add_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exponentnormmode_sub_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exponentnormmode_sub_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_mantissanorm_add_datab	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_mantissanorm_add_result	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_quadrantsum_add_cin	:	STD_LOGIC;
	 SIGNAL  wire_quadrantsum_add_result	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_sft_result	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_cmul_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_lg_negative_quadrant_w19w	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_w_lg_positive_quadrant_w20w	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_circle_w_range7w8w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_input_number_delay_w_range391w392w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_input_number_delay_w_range396w397w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range311w312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range314w315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range317w318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range320w321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range323w324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range326w327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range329w330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range332w333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range335w336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range338w339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range341w342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range344w345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range347w348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range350w351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range353w354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range356w357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range359w360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range362w363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range365w366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range368w369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range371w372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range374w375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range377w378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_negcircle_w_range4w5w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_lg_quadrantselect_w6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_quadrant_w_range17w18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range249w251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range279w281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range282w284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range285w287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range288w290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range291w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range252w254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range255w257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range258w260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range261w263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range264w266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range267w269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range270w272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range273w275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range276w278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_quadrantsign_w57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  circle_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  countnode_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  exponentcheck_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exponentnormmode_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  fixed_sincos_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  fixed_sincosnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  fraction_quadrant_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  indexbit_w :	STD_LOGIC;
	 SIGNAL  indexcheck_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  input_number_delay_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  input_number_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  mantissanormnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  negative_quadrant_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  negcircle_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  one_term_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  overflownode_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  piovertwo_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  positive_quadrant_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  quadrant_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  quadrantselect_w :	STD_LOGIC;
	 SIGNAL  quadrantsign_w :	STD_LOGIC;
	 SIGNAL  radiansnode_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  value_128_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  value_x73_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  zerovec_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_w_circle_w_range7w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_data_range128w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_input_number_delay_w_range391w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_input_number_delay_w_range396w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_negcircle_w_range4w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_quadrant_w_range17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  sinhw_altfp_sincos_cordic_m_e5e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		indexbit	:	IN  STD_LOGIC := '0';
		radians	:	IN  STD_LOGIC_VECTOR(33 DOWNTO 0) := (OTHERS => '0');
		sincos	:	OUT  STD_LOGIC_VECTOR(33 DOWNTO 0);
		sincosbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altfp_sincos_range_b6c
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		circle	:	OUT  STD_LOGIC_VECTOR(35 DOWNTO 0);
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
		negcircle	:	OUT  STD_LOGIC_VECTOR(35 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  sinhw_altpriority_encoder_0c6
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_clshift
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_SHIFTTYPE	:	STRING := "LOGICAL";
		LPM_WIDTH	:	NATURAL;
		LPM_WIDTHDIST	:	NATURAL;
		lpm_type	:	STRING := "lpm_clshift"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		direction	:	IN STD_LOGIC := '0';
		distance	:	IN STD_LOGIC_VECTOR(LPM_WIDTHDIST-1 DOWNTO 0);
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		underflow	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	loop65 : FOR i IN 0 TO 35 GENERATE 
		wire_w_lg_negative_quadrant_w19w(i) <= negative_quadrant_w(i) AND wire_w_lg_w_quadrant_w_range17w18w(0);
	END GENERATE loop65;
	loop66 : FOR i IN 0 TO 35 GENERATE 
		wire_w_lg_positive_quadrant_w20w(i) <= positive_quadrant_w(i) AND wire_w_quadrant_w_range17w(0);
	END GENERATE loop66;
	loop67 : FOR i IN 0 TO 33 GENERATE 
		wire_w_lg_w_circle_w_range7w8w(i) <= wire_w_circle_w_range7w(i) AND wire_w_lg_quadrantselect_w6w(0);
	END GENERATE loop67;
	loop68 : FOR i IN 0 TO 22 GENERATE 
		wire_w_lg_w_input_number_delay_w_range391w392w(i) <= wire_w_input_number_delay_w_range391w(i) AND wire_selectoutputff_w_q_range390w(0);
	END GENERATE loop68;
	loop69 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_input_number_delay_w_range396w397w(i) <= wire_w_input_number_delay_w_range396w(i) AND wire_selectoutputff_w_q_range390w(0);
	END GENERATE loop69;
	wire_w_lg_w_mantissanormnode_w_range311w312w(0) <= wire_w_mantissanormnode_w_range311w(0) AND wire_w_overflownode_w_range309w(0);
	wire_w_lg_w_mantissanormnode_w_range314w315w(0) <= wire_w_mantissanormnode_w_range314w(0) AND wire_w_overflownode_w_range313w(0);
	wire_w_lg_w_mantissanormnode_w_range317w318w(0) <= wire_w_mantissanormnode_w_range317w(0) AND wire_w_overflownode_w_range316w(0);
	wire_w_lg_w_mantissanormnode_w_range320w321w(0) <= wire_w_mantissanormnode_w_range320w(0) AND wire_w_overflownode_w_range319w(0);
	wire_w_lg_w_mantissanormnode_w_range323w324w(0) <= wire_w_mantissanormnode_w_range323w(0) AND wire_w_overflownode_w_range322w(0);
	wire_w_lg_w_mantissanormnode_w_range326w327w(0) <= wire_w_mantissanormnode_w_range326w(0) AND wire_w_overflownode_w_range325w(0);
	wire_w_lg_w_mantissanormnode_w_range329w330w(0) <= wire_w_mantissanormnode_w_range329w(0) AND wire_w_overflownode_w_range328w(0);
	wire_w_lg_w_mantissanormnode_w_range332w333w(0) <= wire_w_mantissanormnode_w_range332w(0) AND wire_w_overflownode_w_range331w(0);
	wire_w_lg_w_mantissanormnode_w_range335w336w(0) <= wire_w_mantissanormnode_w_range335w(0) AND wire_w_overflownode_w_range334w(0);
	wire_w_lg_w_mantissanormnode_w_range338w339w(0) <= wire_w_mantissanormnode_w_range338w(0) AND wire_w_overflownode_w_range337w(0);
	wire_w_lg_w_mantissanormnode_w_range341w342w(0) <= wire_w_mantissanormnode_w_range341w(0) AND wire_w_overflownode_w_range340w(0);
	wire_w_lg_w_mantissanormnode_w_range344w345w(0) <= wire_w_mantissanormnode_w_range344w(0) AND wire_w_overflownode_w_range343w(0);
	wire_w_lg_w_mantissanormnode_w_range347w348w(0) <= wire_w_mantissanormnode_w_range347w(0) AND wire_w_overflownode_w_range346w(0);
	wire_w_lg_w_mantissanormnode_w_range350w351w(0) <= wire_w_mantissanormnode_w_range350w(0) AND wire_w_overflownode_w_range349w(0);
	wire_w_lg_w_mantissanormnode_w_range353w354w(0) <= wire_w_mantissanormnode_w_range353w(0) AND wire_w_overflownode_w_range352w(0);
	wire_w_lg_w_mantissanormnode_w_range356w357w(0) <= wire_w_mantissanormnode_w_range356w(0) AND wire_w_overflownode_w_range355w(0);
	wire_w_lg_w_mantissanormnode_w_range359w360w(0) <= wire_w_mantissanormnode_w_range359w(0) AND wire_w_overflownode_w_range358w(0);
	wire_w_lg_w_mantissanormnode_w_range362w363w(0) <= wire_w_mantissanormnode_w_range362w(0) AND wire_w_overflownode_w_range361w(0);
	wire_w_lg_w_mantissanormnode_w_range365w366w(0) <= wire_w_mantissanormnode_w_range365w(0) AND wire_w_overflownode_w_range364w(0);
	wire_w_lg_w_mantissanormnode_w_range368w369w(0) <= wire_w_mantissanormnode_w_range368w(0) AND wire_w_overflownode_w_range367w(0);
	wire_w_lg_w_mantissanormnode_w_range371w372w(0) <= wire_w_mantissanormnode_w_range371w(0) AND wire_w_overflownode_w_range370w(0);
	wire_w_lg_w_mantissanormnode_w_range374w375w(0) <= wire_w_mantissanormnode_w_range374w(0) AND wire_w_overflownode_w_range373w(0);
	wire_w_lg_w_mantissanormnode_w_range377w378w(0) <= wire_w_mantissanormnode_w_range377w(0) AND wire_w_overflownode_w_range376w(0);
	loop70 : FOR i IN 0 TO 33 GENERATE 
		wire_w_lg_w_negcircle_w_range4w5w(i) <= wire_w_negcircle_w_range4w(i) AND quadrantselect_w;
	END GENERATE loop70;
	wire_w_lg_quadrantselect_w6w(0) <= NOT quadrantselect_w;
	wire_w_lg_w_quadrant_w_range17w18w(0) <= NOT wire_w_quadrant_w_range17w(0);
	wire_w_lg_w_indexcheck_w_range249w251w(0) <= wire_w_indexcheck_w_range249w(0) OR wire_w_radiansnode_w_range248w(0);
	wire_w_lg_w_indexcheck_w_range279w281w(0) <= wire_w_indexcheck_w_range279w(0) OR wire_w_radiansnode_w_range280w(0);
	wire_w_lg_w_indexcheck_w_range282w284w(0) <= wire_w_indexcheck_w_range282w(0) OR wire_w_radiansnode_w_range283w(0);
	wire_w_lg_w_indexcheck_w_range285w287w(0) <= wire_w_indexcheck_w_range285w(0) OR wire_w_radiansnode_w_range286w(0);
	wire_w_lg_w_indexcheck_w_range288w290w(0) <= wire_w_indexcheck_w_range288w(0) OR wire_w_radiansnode_w_range289w(0);
	wire_w_lg_w_indexcheck_w_range291w293w(0) <= wire_w_indexcheck_w_range291w(0) OR wire_w_radiansnode_w_range292w(0);
	wire_w_lg_w_indexcheck_w_range252w254w(0) <= wire_w_indexcheck_w_range252w(0) OR wire_w_radiansnode_w_range253w(0);
	wire_w_lg_w_indexcheck_w_range255w257w(0) <= wire_w_indexcheck_w_range255w(0) OR wire_w_radiansnode_w_range256w(0);
	wire_w_lg_w_indexcheck_w_range258w260w(0) <= wire_w_indexcheck_w_range258w(0) OR wire_w_radiansnode_w_range259w(0);
	wire_w_lg_w_indexcheck_w_range261w263w(0) <= wire_w_indexcheck_w_range261w(0) OR wire_w_radiansnode_w_range262w(0);
	wire_w_lg_w_indexcheck_w_range264w266w(0) <= wire_w_indexcheck_w_range264w(0) OR wire_w_radiansnode_w_range265w(0);
	wire_w_lg_w_indexcheck_w_range267w269w(0) <= wire_w_indexcheck_w_range267w(0) OR wire_w_radiansnode_w_range268w(0);
	wire_w_lg_w_indexcheck_w_range270w272w(0) <= wire_w_indexcheck_w_range270w(0) OR wire_w_radiansnode_w_range271w(0);
	wire_w_lg_w_indexcheck_w_range273w275w(0) <= wire_w_indexcheck_w_range273w(0) OR wire_w_radiansnode_w_range274w(0);
	wire_w_lg_w_indexcheck_w_range276w278w(0) <= wire_w_indexcheck_w_range276w(0) OR wire_w_radiansnode_w_range277w(0);
	wire_w_lg_quadrantsign_w57w(0) <= quadrantsign_w XOR wire_signinff_w_q_range56w(0);
	aclr <= '0';
	circle_w <= wire_crr_fp_range1_circle;
	clk_en <= '1';
	countnode_w <= (NOT wire_clz_q);
	exponentcheck_w <= wire_exponentcheck_sub_result;
	exponentnormmode_w <= wire_exponentnormmode_sub_result;
	fixed_sincos_w <= wire_ccc_cordic_m_sincos;
	fixed_sincosnode_w <= ( fixed_sincos_w & zerovec_w(1 DOWNTO 0));
	fraction_quadrant_w <= (wire_w_lg_positive_quadrant_w20w OR wire_w_lg_negative_quadrant_w19w);
	indexbit_w <= (NOT indexcheck_w(3));
	indexcheck_w <= ( wire_w_lg_w_indexcheck_w_range291w293w & wire_w_lg_w_indexcheck_w_range288w290w & wire_w_lg_w_indexcheck_w_range285w287w & wire_w_lg_w_indexcheck_w_range282w284w & wire_w_lg_w_indexcheck_w_range279w281w & wire_w_lg_w_indexcheck_w_range276w278w & wire_w_lg_w_indexcheck_w_range273w275w & wire_w_lg_w_indexcheck_w_range270w272w & wire_w_lg_w_indexcheck_w_range267w269w & wire_w_lg_w_indexcheck_w_range264w266w & wire_w_lg_w_indexcheck_w_range261w263w & wire_w_lg_w_indexcheck_w_range258w260w & wire_w_lg_w_indexcheck_w_range255w257w & wire_w_lg_w_indexcheck_w_range252w254w & wire_w_lg_w_indexcheck_w_range249w251w & radiansnode_w(32));
	input_number_delay_w <= input_delay_ff_34;
	input_number_w <= data;
	mantissanormnode_w <= wire_sft_result;
	negative_quadrant_w <= (NOT positive_quadrant_w);
	negcircle_w <= wire_crr_fp_range1_negcircle;
	one_term_w <= ( wire_w_lg_w_quadrant_w_range17w18w & zerovec_w(34 DOWNTO 0));
	overflownode_w <= ( wire_w_lg_w_mantissanormnode_w_range377w378w & wire_w_lg_w_mantissanormnode_w_range374w375w & wire_w_lg_w_mantissanormnode_w_range371w372w & wire_w_lg_w_mantissanormnode_w_range368w369w & wire_w_lg_w_mantissanormnode_w_range365w366w & wire_w_lg_w_mantissanormnode_w_range362w363w & wire_w_lg_w_mantissanormnode_w_range359w360w & wire_w_lg_w_mantissanormnode_w_range356w357w & wire_w_lg_w_mantissanormnode_w_range353w354w & wire_w_lg_w_mantissanormnode_w_range350w351w & wire_w_lg_w_mantissanormnode_w_range347w348w & wire_w_lg_w_mantissanormnode_w_range344w345w & wire_w_lg_w_mantissanormnode_w_range341w342w & wire_w_lg_w_mantissanormnode_w_range338w339w & wire_w_lg_w_mantissanormnode_w_range335w336w & wire_w_lg_w_mantissanormnode_w_range332w333w & wire_w_lg_w_mantissanormnode_w_range329w330w & wire_w_lg_w_mantissanormnode_w_range326w327w & wire_w_lg_w_mantissanormnode_w_range323w324w & wire_w_lg_w_mantissanormnode_w_range320w321w & wire_w_lg_w_mantissanormnode_w_range317w318w & wire_w_lg_w_mantissanormnode_w_range314w315w & wire_w_lg_w_mantissanormnode_w_range311w312w & mantissanormnode_w(11));
	piovertwo_w <= "110010010000111111011010101000100010";
	positive_quadrant_w <= ( "0" & quadrant_w & "0");
	quadrant_w <= (wire_w_lg_w_circle_w_range7w8w OR wire_w_lg_w_negcircle_w_range4w5w);
	quadrantselect_w <= circle_w(34);
	quadrantsign_w <= circle_w(35);
	radiansnode_w <= wire_cmul_result;
	result <= ( signoutff & exponentoutff & mantissaoutff);
	value_128_w <= "10000000";
	value_x73_w <= "01110011";
	zerovec_w <= (OTHERS => '0');
	wire_w_circle_w_range7w <= circle_w(33 DOWNTO 0);
	wire_w_data_range128w <= data(30 DOWNTO 23);
	wire_w_indexcheck_w_range249w(0) <= indexcheck_w(0);
	wire_w_indexcheck_w_range279w(0) <= indexcheck_w(10);
	wire_w_indexcheck_w_range282w(0) <= indexcheck_w(11);
	wire_w_indexcheck_w_range285w(0) <= indexcheck_w(12);
	wire_w_indexcheck_w_range288w(0) <= indexcheck_w(13);
	wire_w_indexcheck_w_range291w(0) <= indexcheck_w(14);
	wire_w_indexcheck_w_range252w(0) <= indexcheck_w(1);
	wire_w_indexcheck_w_range255w(0) <= indexcheck_w(2);
	wire_w_indexcheck_w_range258w(0) <= indexcheck_w(3);
	wire_w_indexcheck_w_range261w(0) <= indexcheck_w(4);
	wire_w_indexcheck_w_range264w(0) <= indexcheck_w(5);
	wire_w_indexcheck_w_range267w(0) <= indexcheck_w(6);
	wire_w_indexcheck_w_range270w(0) <= indexcheck_w(7);
	wire_w_indexcheck_w_range273w(0) <= indexcheck_w(8);
	wire_w_indexcheck_w_range276w(0) <= indexcheck_w(9);
	wire_w_input_number_delay_w_range391w <= input_number_delay_w(22 DOWNTO 0);
	wire_w_input_number_delay_w_range396w <= input_number_delay_w(30 DOWNTO 23);
	wire_w_mantissanormnode_w_range311w(0) <= mantissanormnode_w(12);
	wire_w_mantissanormnode_w_range314w(0) <= mantissanormnode_w(13);
	wire_w_mantissanormnode_w_range317w(0) <= mantissanormnode_w(14);
	wire_w_mantissanormnode_w_range320w(0) <= mantissanormnode_w(15);
	wire_w_mantissanormnode_w_range323w(0) <= mantissanormnode_w(16);
	wire_w_mantissanormnode_w_range326w(0) <= mantissanormnode_w(17);
	wire_w_mantissanormnode_w_range329w(0) <= mantissanormnode_w(18);
	wire_w_mantissanormnode_w_range332w(0) <= mantissanormnode_w(19);
	wire_w_mantissanormnode_w_range335w(0) <= mantissanormnode_w(20);
	wire_w_mantissanormnode_w_range338w(0) <= mantissanormnode_w(21);
	wire_w_mantissanormnode_w_range341w(0) <= mantissanormnode_w(22);
	wire_w_mantissanormnode_w_range344w(0) <= mantissanormnode_w(23);
	wire_w_mantissanormnode_w_range347w(0) <= mantissanormnode_w(24);
	wire_w_mantissanormnode_w_range350w(0) <= mantissanormnode_w(25);
	wire_w_mantissanormnode_w_range353w(0) <= mantissanormnode_w(26);
	wire_w_mantissanormnode_w_range356w(0) <= mantissanormnode_w(27);
	wire_w_mantissanormnode_w_range359w(0) <= mantissanormnode_w(28);
	wire_w_mantissanormnode_w_range362w(0) <= mantissanormnode_w(29);
	wire_w_mantissanormnode_w_range365w(0) <= mantissanormnode_w(30);
	wire_w_mantissanormnode_w_range368w(0) <= mantissanormnode_w(31);
	wire_w_mantissanormnode_w_range371w(0) <= mantissanormnode_w(32);
	wire_w_mantissanormnode_w_range374w(0) <= mantissanormnode_w(33);
	wire_w_mantissanormnode_w_range377w(0) <= mantissanormnode_w(34);
	wire_w_negcircle_w_range4w <= negcircle_w(33 DOWNTO 0);
	wire_w_overflownode_w_range309w(0) <= overflownode_w(0);
	wire_w_overflownode_w_range340w(0) <= overflownode_w(10);
	wire_w_overflownode_w_range343w(0) <= overflownode_w(11);
	wire_w_overflownode_w_range346w(0) <= overflownode_w(12);
	wire_w_overflownode_w_range349w(0) <= overflownode_w(13);
	wire_w_overflownode_w_range352w(0) <= overflownode_w(14);
	wire_w_overflownode_w_range355w(0) <= overflownode_w(15);
	wire_w_overflownode_w_range358w(0) <= overflownode_w(16);
	wire_w_overflownode_w_range361w(0) <= overflownode_w(17);
	wire_w_overflownode_w_range364w(0) <= overflownode_w(18);
	wire_w_overflownode_w_range367w(0) <= overflownode_w(19);
	wire_w_overflownode_w_range313w(0) <= overflownode_w(1);
	wire_w_overflownode_w_range370w(0) <= overflownode_w(20);
	wire_w_overflownode_w_range373w(0) <= overflownode_w(21);
	wire_w_overflownode_w_range376w(0) <= overflownode_w(22);
	wire_w_overflownode_w_range316w(0) <= overflownode_w(2);
	wire_w_overflownode_w_range319w(0) <= overflownode_w(3);
	wire_w_overflownode_w_range322w(0) <= overflownode_w(4);
	wire_w_overflownode_w_range325w(0) <= overflownode_w(5);
	wire_w_overflownode_w_range328w(0) <= overflownode_w(6);
	wire_w_overflownode_w_range331w(0) <= overflownode_w(7);
	wire_w_overflownode_w_range334w(0) <= overflownode_w(8);
	wire_w_overflownode_w_range337w(0) <= overflownode_w(9);
	wire_w_quadrant_w_range17w(0) <= quadrant_w(33);
	wire_w_radiansnode_w_range292w(0) <= radiansnode_w(18);
	wire_w_radiansnode_w_range289w(0) <= radiansnode_w(19);
	wire_w_radiansnode_w_range286w(0) <= radiansnode_w(20);
	wire_w_radiansnode_w_range283w(0) <= radiansnode_w(21);
	wire_w_radiansnode_w_range280w(0) <= radiansnode_w(22);
	wire_w_radiansnode_w_range277w(0) <= radiansnode_w(23);
	wire_w_radiansnode_w_range274w(0) <= radiansnode_w(24);
	wire_w_radiansnode_w_range271w(0) <= radiansnode_w(25);
	wire_w_radiansnode_w_range268w(0) <= radiansnode_w(26);
	wire_w_radiansnode_w_range265w(0) <= radiansnode_w(27);
	wire_w_radiansnode_w_range262w(0) <= radiansnode_w(28);
	wire_w_radiansnode_w_range259w(0) <= radiansnode_w(29);
	wire_w_radiansnode_w_range256w(0) <= radiansnode_w(30);
	wire_w_radiansnode_w_range253w(0) <= radiansnode_w(31);
	wire_w_radiansnode_w_range248w(0) <= radiansnode_w(32);
	ccc_cordic_m :  sinhw_altfp_sincos_cordic_m_e5e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		indexbit => indexbit_w,
		radians => radiansnode_w,
		sincos => wire_ccc_cordic_m_sincos,
		sincosbit => select_sincosff(3)
	  );
	crr_fp_range1 :  sinhw_altfp_sincos_range_b6c
	  PORT MAP ( 
		aclr => aclr,
		circle => wire_crr_fp_range1_circle,
		clken => clk_en,
		clock => clock,
		data => data,
		negcircle => wire_crr_fp_range1_negcircle
	  );
	wire_clz_data <= ( fixed_sincosnode_w & "1111111111111111111111111111");
	clz :  sinhw_altpriority_encoder_0c6
	  PORT MAP ( 
		data => wire_clz_data,
		q => wire_clz_q
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN countff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN countff <= countnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponentinff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponentinff <= wire_w_data_range128w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponentnormff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponentnormff <= wire_exponentnorm_add_result;
			END IF;
		END IF;
	END PROCESS;
	loop71 : FOR i IN 0 TO 7 GENERATE 
		wire_exponentnormff_w_lg_q398w(i) <= exponentnormff(i) AND wire_selectoutputff_w_lg_w_q_range390w393w(0);
	END GENERATE loop71;
	loop72 : FOR i IN 0 TO 7 GENERATE 
		wire_exponentnormff_w_lg_w_lg_q398w399w(i) <= wire_exponentnormff_w_lg_q398w(i) OR wire_w_lg_w_input_number_delay_w_range396w397w(i);
	END GENERATE loop72;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponentoutff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponentoutff <= wire_exponentnormff_w_lg_w_lg_q398w399w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN fixed_sincosff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN fixed_sincosff <= fixed_sincosnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_0 <= input_number_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_1 <= input_delay_ff_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_10 <= input_delay_ff_9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_11 <= input_delay_ff_10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_12 <= input_delay_ff_11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_13 <= input_delay_ff_12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_14 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_14 <= input_delay_ff_13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_15 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_15 <= input_delay_ff_14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_16 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_16 <= input_delay_ff_15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_17 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_17 <= input_delay_ff_16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_18 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_18 <= input_delay_ff_17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_19 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_19 <= input_delay_ff_18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_2 <= input_delay_ff_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_20 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_20 <= input_delay_ff_19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_21 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_21 <= input_delay_ff_20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_22 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_22 <= input_delay_ff_21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_23 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_23 <= input_delay_ff_22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_24 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_24 <= input_delay_ff_23;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_25 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_25 <= input_delay_ff_24;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_26 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_26 <= input_delay_ff_25;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_27 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_27 <= input_delay_ff_26;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_28 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_28 <= input_delay_ff_27;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_29 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_29 <= input_delay_ff_28;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_3 <= input_delay_ff_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_30 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_30 <= input_delay_ff_29;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_31 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_31 <= input_delay_ff_30;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_32 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_32 <= input_delay_ff_31;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_33 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_33 <= input_delay_ff_32;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_34 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_34 <= input_delay_ff_33;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_4 <= input_delay_ff_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_5 <= input_delay_ff_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_6 <= input_delay_ff_5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_7 <= input_delay_ff_6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_8 <= input_delay_ff_7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN input_delay_ff_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN input_delay_ff_9 <= input_delay_ff_8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissanormff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissanormff <= wire_mantissanorm_add_result;
			END IF;
		END IF;
	END PROCESS;
	loop73 : FOR i IN 0 TO 22 GENERATE 
		wire_mantissanormff_w_lg_q394w(i) <= mantissanormff(i) AND wire_selectoutputff_w_lg_w_q_range390w393w(0);
	END GENERATE loop73;
	loop74 : FOR i IN 0 TO 22 GENERATE 
		wire_mantissanormff_w_lg_w_lg_q394w395w(i) <= wire_mantissanormff_w_lg_q394w(i) OR wire_w_lg_w_input_number_delay_w_range391w392w(i);
	END GENERATE loop74;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissaoutff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissaoutff <= wire_mantissanormff_w_lg_w_lg_q394w395w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN quadrant_sumff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN quadrant_sumff <= wire_quadrantsum_add_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN select_sincosff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN select_sincosff <= ( select_sincosff(2 DOWNTO 0) & quadrant_w(33));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN selectoutputff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN selectoutputff <= ( selectoutputff(32 DOWNTO 0) & exponentcheck_w(8));
			END IF;
		END IF;
	END PROCESS;
	wire_selectoutputff_w_lg_w_q_range390w393w(0) <= NOT wire_selectoutputff_w_q_range390w(0);
	wire_selectoutputff_w_q_range390w(0) <= selectoutputff(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN signcalcff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN signcalcff <= ( signcalcff(22 DOWNTO 0) & wire_w_lg_quadrantsign_w57w);
			END IF;
		END IF;
	END PROCESS;
	wire_signcalcff_w_lg_w_q_range402w403w(0) <= wire_signcalcff_w_q_range402w(0) AND wire_selectoutputff_w_lg_w_q_range390w393w(0);
	wire_signcalcff_w_q_range402w(0) <= signcalcff(23);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN signinff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN signinff <= ( signinff(9 DOWNTO 0) & data(31));
			END IF;
		END IF;
	END PROCESS;
	wire_signinff_w_q_range56w(0) <= signinff(10);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN signoutff <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN signoutff <= (wire_signcalcff_w_lg_w_q_range402w403w(0) OR (input_number_delay_w(31) AND selectoutputff(33)));
			END IF;
		END IF;
	END PROCESS;
	wire_exponentcheck_sub_dataa <= ( "0" & exponentinff);
	wire_exponentcheck_sub_datab <= ( "0" & value_x73_w);
	exponentcheck_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => wire_exponentcheck_sub_dataa,
		datab => wire_exponentcheck_sub_datab,
		result => wire_exponentcheck_sub_result
	  );
	wire_exponentnorm_add_datab <= ( "0000000" & overflownode_w(23));
	exponentnorm_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		dataa => exponentnormmode_w(7 DOWNTO 0),
		datab => wire_exponentnorm_add_datab,
		result => wire_exponentnorm_add_result
	  );
	wire_exponentnormmode_sub_datab <= ( "00" & countff);
	exponentnormmode_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		dataa => value_128_w,
		datab => wire_exponentnormmode_sub_datab,
		result => wire_exponentnormmode_sub_result
	  );
	wire_mantissanorm_add_datab <= ( "0000000000000000000000" & mantissanormnode_w(11));
	mantissanorm_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 23
	  )
	  PORT MAP ( 
		dataa => mantissanormnode_w(34 DOWNTO 12),
		datab => wire_mantissanorm_add_datab,
		result => wire_mantissanorm_add_result
	  );
	wire_quadrantsum_add_cin <= wire_w_lg_w_quadrant_w_range17w18w(0);
	quadrantsum_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 36
	  )
	  PORT MAP ( 
		cin => wire_quadrantsum_add_cin,
		dataa => one_term_w,
		datab => fraction_quadrant_w,
		result => wire_quadrantsum_add_result
	  );
	sft :  lpm_clshift
	  GENERIC MAP (
		LPM_WIDTH => 36,
		LPM_WIDTHDIST => 6
	  )
	  PORT MAP ( 
		data => fixed_sincosff,
		direction => wire_gnd,
		distance => countff,
		result => wire_sft_result
	  );
	cmul :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 36,
		LPM_WIDTHB => 36,
		LPM_WIDTHP => 34
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => quadrant_sumff,
		datab => piovertwo_w,
		result => wire_cmul_result
	  );

 END RTL; --sinhw_altfp_sincos_47e
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY sinhw IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END sinhw;


ARCHITECTURE RTL OF sinhw IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT sinhw_altfp_sincos_47e
	PORT (
			clock	: IN STD_LOGIC ;
			data	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	sinhw_altfp_sincos_47e_component : sinhw_altfp_sincos_47e
	PORT MAP (
		clock => clock,
		data => data,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: FPM_FORMAT NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: OPERATION STRING "SIN"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "36"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data 0 0 32 0 INPUT NODEFVAL "data[31..0]"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data 0 0 32 0 data 0 0 32 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL sinhw.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sinhw.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sinhw.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sinhw.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL sinhw_inst.vhd FALSE
