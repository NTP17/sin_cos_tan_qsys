-- firmware.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity firmware is
	port (
		clk_clk          : in  std_logic                     := '0'; --     clk.clk
		cos_out_readdata : out std_logic_vector(31 downto 0);        -- cos_out.readdata
		pio_out_export   : out std_logic_vector(31 downto 0);        -- pio_out.export
		reset_reset_n    : in  std_logic                     := '0'; --   reset.reset_n
		sin_out_readdata : out std_logic_vector(31 downto 0);        -- sin_out.readdata
		tan_out_readdata : out std_logic_vector(31 downto 0)         -- tan_out.readdata
	);
end entity firmware;

architecture rtl of firmware is
	component hwcos is
		port (
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			chipselect : in  std_logic                     := 'X';             -- chipselect
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			clock      : in  std_logic                     := 'X';             -- clk
			conduit    : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component hwcos;

	component firmware_CPU is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(19 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(19 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component firmware_CPU;

	component firmware_MEMORY is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component firmware_MEMORY;

	component firmware_PIO is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component firmware_PIO;

	component hwsin is
		port (
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			chipselect : in  std_logic                     := 'X';             -- chipselect
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			conduit    : out std_logic_vector(31 downto 0);                    -- readdata
			clock      : in  std_logic                     := 'X'              -- clk
		);
	end component hwsin;

	component hwtan is
		port (
			read       : in  std_logic                     := 'X';             -- read
			write      : in  std_logic                     := 'X';             -- write
			chipselect : in  std_logic                     := 'X';             -- chipselect
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			clock      : in  std_logic                     := 'X';             -- clk
			conduit    : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component hwtan;

	component firmware_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component firmware_jtag_uart_0;

	component firmware_mm_interconnect_0 is
		port (
			clk_0_clk_clk                             : in  std_logic                     := 'X';             -- clk
			CPU_reset_reset_bridge_in_reset_reset     : in  std_logic                     := 'X';             -- reset
			CPU_data_master_address                   : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			CPU_data_master_waitrequest               : out std_logic;                                        -- waitrequest
			CPU_data_master_byteenable                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			CPU_data_master_read                      : in  std_logic                     := 'X';             -- read
			CPU_data_master_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_data_master_readdatavalid             : out std_logic;                                        -- readdatavalid
			CPU_data_master_write                     : in  std_logic                     := 'X';             -- write
			CPU_data_master_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_data_master_debugaccess               : in  std_logic                     := 'X';             -- debugaccess
			CPU_instruction_master_address            : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			CPU_instruction_master_waitrequest        : out std_logic;                                        -- waitrequest
			CPU_instruction_master_read               : in  std_logic                     := 'X';             -- read
			CPU_instruction_master_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_instruction_master_readdatavalid      : out std_logic;                                        -- readdatavalid
			COS_HW_avalon_slave_0_write               : out std_logic;                                        -- write
			COS_HW_avalon_slave_0_read                : out std_logic;                                        -- read
			COS_HW_avalon_slave_0_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			COS_HW_avalon_slave_0_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			COS_HW_avalon_slave_0_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			COS_HW_avalon_slave_0_chipselect          : out std_logic;                                        -- chipselect
			CPU_debug_mem_slave_address               : out std_logic_vector(8 downto 0);                     -- address
			CPU_debug_mem_slave_write                 : out std_logic;                                        -- write
			CPU_debug_mem_slave_read                  : out std_logic;                                        -- read
			CPU_debug_mem_slave_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_debug_mem_slave_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_debug_mem_slave_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			CPU_debug_mem_slave_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			CPU_debug_mem_slave_debugaccess           : out std_logic;                                        -- debugaccess
			jtag_uart_0_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			MEMORY_s1_address                         : out std_logic_vector(15 downto 0);                    -- address
			MEMORY_s1_write                           : out std_logic;                                        -- write
			MEMORY_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			MEMORY_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			MEMORY_s1_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			MEMORY_s1_chipselect                      : out std_logic;                                        -- chipselect
			MEMORY_s1_clken                           : out std_logic;                                        -- clken
			PIO_s1_address                            : out std_logic_vector(1 downto 0);                     -- address
			PIO_s1_write                              : out std_logic;                                        -- write
			PIO_s1_readdata                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PIO_s1_writedata                          : out std_logic_vector(31 downto 0);                    -- writedata
			PIO_s1_chipselect                         : out std_logic;                                        -- chipselect
			SIN_HW_avalon_slave_0_write               : out std_logic;                                        -- write
			SIN_HW_avalon_slave_0_read                : out std_logic;                                        -- read
			SIN_HW_avalon_slave_0_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SIN_HW_avalon_slave_0_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			SIN_HW_avalon_slave_0_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			SIN_HW_avalon_slave_0_chipselect          : out std_logic;                                        -- chipselect
			TAN_HW_avalon_slave_0_write               : out std_logic;                                        -- write
			TAN_HW_avalon_slave_0_read                : out std_logic;                                        -- read
			TAN_HW_avalon_slave_0_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TAN_HW_avalon_slave_0_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			TAN_HW_avalon_slave_0_byteenable          : out std_logic_vector(3 downto 0);                     -- byteenable
			TAN_HW_avalon_slave_0_chipselect          : out std_logic                                         -- chipselect
		);
	end component firmware_mm_interconnect_0;

	component firmware_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component firmware_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal cpu_data_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	signal cpu_data_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	signal cpu_data_master_debugaccess                                     : std_logic;                     -- CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	signal cpu_data_master_address                                         : std_logic_vector(19 downto 0); -- CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	signal cpu_data_master_byteenable                                      : std_logic_vector(3 downto 0);  -- CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	signal cpu_data_master_read                                            : std_logic;                     -- CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	signal cpu_data_master_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:CPU_data_master_readdatavalid -> CPU:d_readdatavalid
	signal cpu_data_master_write                                           : std_logic;                     -- CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	signal cpu_data_master_writedata                                       : std_logic_vector(31 downto 0); -- CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	signal cpu_instruction_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	signal cpu_instruction_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	signal cpu_instruction_master_address                                  : std_logic_vector(19 downto 0); -- CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	signal cpu_instruction_master_read                                     : std_logic;                     -- CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	signal cpu_instruction_master_readdatavalid                            : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_readdatavalid -> CPU:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_sin_hw_avalon_slave_0_chipselect              : std_logic;                     -- mm_interconnect_0:SIN_HW_avalon_slave_0_chipselect -> SIN_HW:chipselect
	signal mm_interconnect_0_sin_hw_avalon_slave_0_readdata                : std_logic_vector(31 downto 0); -- SIN_HW:readdata -> mm_interconnect_0:SIN_HW_avalon_slave_0_readdata
	signal mm_interconnect_0_sin_hw_avalon_slave_0_read                    : std_logic;                     -- mm_interconnect_0:SIN_HW_avalon_slave_0_read -> SIN_HW:read
	signal mm_interconnect_0_sin_hw_avalon_slave_0_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:SIN_HW_avalon_slave_0_byteenable -> SIN_HW:byteenable
	signal mm_interconnect_0_sin_hw_avalon_slave_0_write                   : std_logic;                     -- mm_interconnect_0:SIN_HW_avalon_slave_0_write -> SIN_HW:write
	signal mm_interconnect_0_sin_hw_avalon_slave_0_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:SIN_HW_avalon_slave_0_writedata -> SIN_HW:writedata
	signal mm_interconnect_0_cos_hw_avalon_slave_0_chipselect              : std_logic;                     -- mm_interconnect_0:COS_HW_avalon_slave_0_chipselect -> COS_HW:chipselect
	signal mm_interconnect_0_cos_hw_avalon_slave_0_readdata                : std_logic_vector(31 downto 0); -- COS_HW:readdata -> mm_interconnect_0:COS_HW_avalon_slave_0_readdata
	signal mm_interconnect_0_cos_hw_avalon_slave_0_read                    : std_logic;                     -- mm_interconnect_0:COS_HW_avalon_slave_0_read -> COS_HW:read
	signal mm_interconnect_0_cos_hw_avalon_slave_0_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:COS_HW_avalon_slave_0_byteenable -> COS_HW:byteenable
	signal mm_interconnect_0_cos_hw_avalon_slave_0_write                   : std_logic;                     -- mm_interconnect_0:COS_HW_avalon_slave_0_write -> COS_HW:write
	signal mm_interconnect_0_cos_hw_avalon_slave_0_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:COS_HW_avalon_slave_0_writedata -> COS_HW:writedata
	signal mm_interconnect_0_tan_hw_avalon_slave_0_chipselect              : std_logic;                     -- mm_interconnect_0:TAN_HW_avalon_slave_0_chipselect -> TAN_HW:chipselect
	signal mm_interconnect_0_tan_hw_avalon_slave_0_readdata                : std_logic_vector(31 downto 0); -- TAN_HW:readdata -> mm_interconnect_0:TAN_HW_avalon_slave_0_readdata
	signal mm_interconnect_0_tan_hw_avalon_slave_0_read                    : std_logic;                     -- mm_interconnect_0:TAN_HW_avalon_slave_0_read -> TAN_HW:read
	signal mm_interconnect_0_tan_hw_avalon_slave_0_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:TAN_HW_avalon_slave_0_byteenable -> TAN_HW:byteenable
	signal mm_interconnect_0_tan_hw_avalon_slave_0_write                   : std_logic;                     -- mm_interconnect_0:TAN_HW_avalon_slave_0_write -> TAN_HW:write
	signal mm_interconnect_0_tan_hw_avalon_slave_0_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:TAN_HW_avalon_slave_0_writedata -> TAN_HW:writedata
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                  : std_logic_vector(31 downto 0); -- CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest               : std_logic;                     -- CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess               : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                   : std_logic_vector(8 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                      : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                     : std_logic;                     -- mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	signal mm_interconnect_0_memory_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:MEMORY_s1_chipselect -> MEMORY:chipselect
	signal mm_interconnect_0_memory_s1_readdata                            : std_logic_vector(31 downto 0); -- MEMORY:readdata -> mm_interconnect_0:MEMORY_s1_readdata
	signal mm_interconnect_0_memory_s1_address                             : std_logic_vector(15 downto 0); -- mm_interconnect_0:MEMORY_s1_address -> MEMORY:address
	signal mm_interconnect_0_memory_s1_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:MEMORY_s1_byteenable -> MEMORY:byteenable
	signal mm_interconnect_0_memory_s1_write                               : std_logic;                     -- mm_interconnect_0:MEMORY_s1_write -> MEMORY:write
	signal mm_interconnect_0_memory_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:MEMORY_s1_writedata -> MEMORY:writedata
	signal mm_interconnect_0_memory_s1_clken                               : std_logic;                     -- mm_interconnect_0:MEMORY_s1_clken -> MEMORY:clken
	signal mm_interconnect_0_pio_s1_chipselect                             : std_logic;                     -- mm_interconnect_0:PIO_s1_chipselect -> PIO:chipselect
	signal mm_interconnect_0_pio_s1_readdata                               : std_logic_vector(31 downto 0); -- PIO:readdata -> mm_interconnect_0:PIO_s1_readdata
	signal mm_interconnect_0_pio_s1_address                                : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PIO_s1_address -> PIO:address
	signal mm_interconnect_0_pio_s1_write                                  : std_logic;                     -- mm_interconnect_0:PIO_s1_write -> mm_interconnect_0_pio_s1_write:in
	signal mm_interconnect_0_pio_s1_writedata                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:PIO_s1_writedata -> PIO:writedata
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal cpu_irq_irq                                                     : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> CPU:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [MEMORY:reset, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [CPU:reset_req, MEMORY:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_pio_s1_write_ports_inv                        : std_logic;                     -- mm_interconnect_0_pio_s1_write:inv -> PIO:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [COS_HW:reset_n, CPU:reset_n, PIO:reset_n, SIN_HW:reset_n, TAN_HW:reset_n, jtag_uart_0:rst_n]

begin

	cos_hw : component hwcos
		port map (
			read       => mm_interconnect_0_cos_hw_avalon_slave_0_read,       -- avalon_slave_0.read
			write      => mm_interconnect_0_cos_hw_avalon_slave_0_write,      --               .write
			chipselect => mm_interconnect_0_cos_hw_avalon_slave_0_chipselect, --               .chipselect
			byteenable => mm_interconnect_0_cos_hw_avalon_slave_0_byteenable, --               .byteenable
			writedata  => mm_interconnect_0_cos_hw_avalon_slave_0_writedata,  --               .writedata
			readdata   => mm_interconnect_0_cos_hw_avalon_slave_0_readdata,   --               .readdata
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --          reset.reset_n
			clock      => clk_clk,                                            --          clock.clk
			conduit    => cos_out_readdata                                    --    conduit_end.readdata
		);

	cpu : component firmware_CPU
		port map (
			clk                                 => clk_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                              --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	memory : component firmware_MEMORY
		port map (
			clk        => clk_clk,                                --   clk1.clk
			address    => mm_interconnect_0_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,         -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,     --       .reset_req
			freeze     => '0'                                     -- (terminated)
		);

	pio : component firmware_PIO
		port map (
			clk        => clk_clk,                                  --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_s1_readdata,        --                    .readdata
			out_port   => pio_out_export                            -- external_connection.export
		);

	sin_hw : component hwsin
		port map (
			read       => mm_interconnect_0_sin_hw_avalon_slave_0_read,       -- avalon_slave_0.read
			write      => mm_interconnect_0_sin_hw_avalon_slave_0_write,      --               .write
			chipselect => mm_interconnect_0_sin_hw_avalon_slave_0_chipselect, --               .chipselect
			byteenable => mm_interconnect_0_sin_hw_avalon_slave_0_byteenable, --               .byteenable
			writedata  => mm_interconnect_0_sin_hw_avalon_slave_0_writedata,  --               .writedata
			readdata   => mm_interconnect_0_sin_hw_avalon_slave_0_readdata,   --               .readdata
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --          reset.reset_n
			conduit    => sin_out_readdata,                                   --    conduit_end.readdata
			clock      => clk_clk                                             --          clock.clk
		);

	tan_hw : component hwtan
		port map (
			read       => mm_interconnect_0_tan_hw_avalon_slave_0_read,       -- avalon_slave_0.read
			write      => mm_interconnect_0_tan_hw_avalon_slave_0_write,      --               .write
			chipselect => mm_interconnect_0_tan_hw_avalon_slave_0_chipselect, --               .chipselect
			byteenable => mm_interconnect_0_tan_hw_avalon_slave_0_byteenable, --               .byteenable
			writedata  => mm_interconnect_0_tan_hw_avalon_slave_0_writedata,  --               .writedata
			readdata   => mm_interconnect_0_tan_hw_avalon_slave_0_readdata,   --               .readdata
			reset_n    => rst_controller_reset_out_reset_ports_inv,           --          reset.reset_n
			clock      => clk_clk,                                            --          clock.clk
			conduit    => tan_out_readdata                                    --    conduit_end.readdata
		);

	jtag_uart_0 : component firmware_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	mm_interconnect_0 : component firmware_mm_interconnect_0
		port map (
			clk_0_clk_clk                             => clk_clk,                                                     --                       clk_0_clk.clk
			CPU_reset_reset_bridge_in_reset_reset     => rst_controller_reset_out_reset,                              -- CPU_reset_reset_bridge_in_reset.reset
			CPU_data_master_address                   => cpu_data_master_address,                                     --                 CPU_data_master.address
			CPU_data_master_waitrequest               => cpu_data_master_waitrequest,                                 --                                .waitrequest
			CPU_data_master_byteenable                => cpu_data_master_byteenable,                                  --                                .byteenable
			CPU_data_master_read                      => cpu_data_master_read,                                        --                                .read
			CPU_data_master_readdata                  => cpu_data_master_readdata,                                    --                                .readdata
			CPU_data_master_readdatavalid             => cpu_data_master_readdatavalid,                               --                                .readdatavalid
			CPU_data_master_write                     => cpu_data_master_write,                                       --                                .write
			CPU_data_master_writedata                 => cpu_data_master_writedata,                                   --                                .writedata
			CPU_data_master_debugaccess               => cpu_data_master_debugaccess,                                 --                                .debugaccess
			CPU_instruction_master_address            => cpu_instruction_master_address,                              --          CPU_instruction_master.address
			CPU_instruction_master_waitrequest        => cpu_instruction_master_waitrequest,                          --                                .waitrequest
			CPU_instruction_master_read               => cpu_instruction_master_read,                                 --                                .read
			CPU_instruction_master_readdata           => cpu_instruction_master_readdata,                             --                                .readdata
			CPU_instruction_master_readdatavalid      => cpu_instruction_master_readdatavalid,                        --                                .readdatavalid
			COS_HW_avalon_slave_0_write               => mm_interconnect_0_cos_hw_avalon_slave_0_write,               --           COS_HW_avalon_slave_0.write
			COS_HW_avalon_slave_0_read                => mm_interconnect_0_cos_hw_avalon_slave_0_read,                --                                .read
			COS_HW_avalon_slave_0_readdata            => mm_interconnect_0_cos_hw_avalon_slave_0_readdata,            --                                .readdata
			COS_HW_avalon_slave_0_writedata           => mm_interconnect_0_cos_hw_avalon_slave_0_writedata,           --                                .writedata
			COS_HW_avalon_slave_0_byteenable          => mm_interconnect_0_cos_hw_avalon_slave_0_byteenable,          --                                .byteenable
			COS_HW_avalon_slave_0_chipselect          => mm_interconnect_0_cos_hw_avalon_slave_0_chipselect,          --                                .chipselect
			CPU_debug_mem_slave_address               => mm_interconnect_0_cpu_debug_mem_slave_address,               --             CPU_debug_mem_slave.address
			CPU_debug_mem_slave_write                 => mm_interconnect_0_cpu_debug_mem_slave_write,                 --                                .write
			CPU_debug_mem_slave_read                  => mm_interconnect_0_cpu_debug_mem_slave_read,                  --                                .read
			CPU_debug_mem_slave_readdata              => mm_interconnect_0_cpu_debug_mem_slave_readdata,              --                                .readdata
			CPU_debug_mem_slave_writedata             => mm_interconnect_0_cpu_debug_mem_slave_writedata,             --                                .writedata
			CPU_debug_mem_slave_byteenable            => mm_interconnect_0_cpu_debug_mem_slave_byteenable,            --                                .byteenable
			CPU_debug_mem_slave_waitrequest           => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,           --                                .waitrequest
			CPU_debug_mem_slave_debugaccess           => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,           --                                .debugaccess
			jtag_uart_0_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --   jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                .write
			jtag_uart_0_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                .read
			jtag_uart_0_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                .readdata
			jtag_uart_0_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                .chipselect
			MEMORY_s1_address                         => mm_interconnect_0_memory_s1_address,                         --                       MEMORY_s1.address
			MEMORY_s1_write                           => mm_interconnect_0_memory_s1_write,                           --                                .write
			MEMORY_s1_readdata                        => mm_interconnect_0_memory_s1_readdata,                        --                                .readdata
			MEMORY_s1_writedata                       => mm_interconnect_0_memory_s1_writedata,                       --                                .writedata
			MEMORY_s1_byteenable                      => mm_interconnect_0_memory_s1_byteenable,                      --                                .byteenable
			MEMORY_s1_chipselect                      => mm_interconnect_0_memory_s1_chipselect,                      --                                .chipselect
			MEMORY_s1_clken                           => mm_interconnect_0_memory_s1_clken,                           --                                .clken
			PIO_s1_address                            => mm_interconnect_0_pio_s1_address,                            --                          PIO_s1.address
			PIO_s1_write                              => mm_interconnect_0_pio_s1_write,                              --                                .write
			PIO_s1_readdata                           => mm_interconnect_0_pio_s1_readdata,                           --                                .readdata
			PIO_s1_writedata                          => mm_interconnect_0_pio_s1_writedata,                          --                                .writedata
			PIO_s1_chipselect                         => mm_interconnect_0_pio_s1_chipselect,                         --                                .chipselect
			SIN_HW_avalon_slave_0_write               => mm_interconnect_0_sin_hw_avalon_slave_0_write,               --           SIN_HW_avalon_slave_0.write
			SIN_HW_avalon_slave_0_read                => mm_interconnect_0_sin_hw_avalon_slave_0_read,                --                                .read
			SIN_HW_avalon_slave_0_readdata            => mm_interconnect_0_sin_hw_avalon_slave_0_readdata,            --                                .readdata
			SIN_HW_avalon_slave_0_writedata           => mm_interconnect_0_sin_hw_avalon_slave_0_writedata,           --                                .writedata
			SIN_HW_avalon_slave_0_byteenable          => mm_interconnect_0_sin_hw_avalon_slave_0_byteenable,          --                                .byteenable
			SIN_HW_avalon_slave_0_chipselect          => mm_interconnect_0_sin_hw_avalon_slave_0_chipselect,          --                                .chipselect
			TAN_HW_avalon_slave_0_write               => mm_interconnect_0_tan_hw_avalon_slave_0_write,               --           TAN_HW_avalon_slave_0.write
			TAN_HW_avalon_slave_0_read                => mm_interconnect_0_tan_hw_avalon_slave_0_read,                --                                .read
			TAN_HW_avalon_slave_0_readdata            => mm_interconnect_0_tan_hw_avalon_slave_0_readdata,            --                                .readdata
			TAN_HW_avalon_slave_0_writedata           => mm_interconnect_0_tan_hw_avalon_slave_0_writedata,           --                                .writedata
			TAN_HW_avalon_slave_0_byteenable          => mm_interconnect_0_tan_hw_avalon_slave_0_byteenable,          --                                .byteenable
			TAN_HW_avalon_slave_0_chipselect          => mm_interconnect_0_tan_hw_avalon_slave_0_chipselect           --                                .chipselect
		);

	irq_mapper : component firmware_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_pio_s1_write_ports_inv <= not mm_interconnect_0_pio_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of firmware
