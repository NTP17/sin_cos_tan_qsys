-- megafunction wizard: %ALTFP_SINCOS%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altfp_sincos 

-- ============================================================
-- File Name: coshw.vhd
-- Megafunction Name(s):
-- 			altfp_sincos
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


--altfp_sincos CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" OPERATION="COS" PIPELINE=35 ROUNDING="TO_NEAREST" WIDTH_EXP=8 WIDTH_MAN=23 clock data result
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END


--altfp_sincos_cordic_m CBX_AUTO_BLACKBOX="ALL" DEPTH=18 DEVICE_FAMILY="Cyclone V" INDEXPOINT=3 WIDTH=32 aclr clken clock indexbit radians sincos sincosbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=0 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_35b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_35b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_35b IS

	 SIGNAL  wire_cata_0_cordic_atan_w_lg_w_lg_indexbit10156w10157w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_0_cordic_atan_w_lg_indexbit10154w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_0_cordic_atan_w_lg_indexbit10156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_0_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_3_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_0_cordic_atan_w_valuenode_0_w_range10155w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_0_cordic_atan_w_valuenode_3_w_range10153w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop0 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_0_cordic_atan_w_lg_w_lg_indexbit10156w10157w(i) <= wire_cata_0_cordic_atan_w_lg_indexbit10156w(0) AND wire_cata_0_cordic_atan_w_valuenode_0_w_range10155w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_0_cordic_atan_w_lg_indexbit10154w(i) <= indexbit AND wire_cata_0_cordic_atan_w_valuenode_3_w_range10153w(i);
	END GENERATE loop1;
	wire_cata_0_cordic_atan_w_lg_indexbit10156w(0) <= NOT indexbit;
	arctan <= (wire_cata_0_cordic_atan_w_lg_w_lg_indexbit10156w10157w OR wire_cata_0_cordic_atan_w_lg_indexbit10154w);
	valuenode_0_w <= "001100100100001111110110101010001000100001011010";
	valuenode_3_w <= "000001111111010101101110101001101010101100001100";
	wire_cata_0_cordic_atan_w_valuenode_0_w_range10155w <= valuenode_0_w(47 DOWNTO 16);
	wire_cata_0_cordic_atan_w_valuenode_3_w_range10153w <= valuenode_3_w(44 DOWNTO 13);

 END RTL; --coshw_altfp_sincos_cordic_atan_35b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=10 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_k6b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_k6b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_k6b IS

	 SIGNAL  wire_cata_10_cordic_atan_w_lg_w_lg_indexbit10162w10163w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_w_lg_indexbit10160w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_w_lg_indexbit10162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_10_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_13_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_w_valuenode_10_w_range10161w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_w_valuenode_13_w_range10159w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop2 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_10_cordic_atan_w_lg_w_lg_indexbit10162w10163w(i) <= wire_cata_10_cordic_atan_w_lg_indexbit10162w(0) AND wire_cata_10_cordic_atan_w_valuenode_10_w_range10161w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_10_cordic_atan_w_lg_indexbit10160w(i) <= indexbit AND wire_cata_10_cordic_atan_w_valuenode_13_w_range10159w(i);
	END GENERATE loop3;
	wire_cata_10_cordic_atan_w_lg_indexbit10162w(0) <= NOT indexbit;
	arctan <= (wire_cata_10_cordic_atan_w_lg_w_lg_indexbit10162w10163w OR wire_cata_10_cordic_atan_w_lg_indexbit10160w);
	valuenode_10_w <= "000000000000111111111111111111111010101010101011";
	valuenode_13_w <= "000000000000000111111111111111111111111111010101";
	wire_cata_10_cordic_atan_w_valuenode_10_w_range10161w <= valuenode_10_w(47 DOWNTO 16);
	wire_cata_10_cordic_atan_w_valuenode_13_w_range10159w <= valuenode_13_w(44 DOWNTO 13);

 END RTL; --coshw_altfp_sincos_cordic_atan_k6b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=11 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_l6b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_l6b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_l6b IS

	 SIGNAL  wire_cata_11_cordic_atan_w_lg_w_lg_indexbit10168w10169w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_w_lg_indexbit10166w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_w_lg_indexbit10168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_11_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_14_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_w_valuenode_11_w_range10167w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_w_valuenode_14_w_range10165w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop4 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_11_cordic_atan_w_lg_w_lg_indexbit10168w10169w(i) <= wire_cata_11_cordic_atan_w_lg_indexbit10168w(0) AND wire_cata_11_cordic_atan_w_valuenode_11_w_range10167w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_11_cordic_atan_w_lg_indexbit10166w(i) <= indexbit AND wire_cata_11_cordic_atan_w_valuenode_14_w_range10165w(i);
	END GENERATE loop5;
	wire_cata_11_cordic_atan_w_lg_indexbit10168w(0) <= NOT indexbit;
	arctan <= (wire_cata_11_cordic_atan_w_lg_w_lg_indexbit10168w10169w OR wire_cata_11_cordic_atan_w_lg_indexbit10166w);
	valuenode_11_w <= "000000000000011111111111111111111111010101010101";
	valuenode_14_w <= "000000000000000011111111111111111111111111111011";
	wire_cata_11_cordic_atan_w_valuenode_11_w_range10167w <= valuenode_11_w(47 DOWNTO 16);
	wire_cata_11_cordic_atan_w_valuenode_14_w_range10165w <= valuenode_14_w(44 DOWNTO 13);

 END RTL; --coshw_altfp_sincos_cordic_atan_l6b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=12 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_m6b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_m6b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_m6b IS

	 SIGNAL  wire_cata_12_cordic_atan_w_lg_w_lg_indexbit10174w10175w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_w_lg_indexbit10172w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_w_lg_indexbit10174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_12_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_15_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_w_valuenode_12_w_range10173w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_w_valuenode_15_w_range10171w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop6 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_12_cordic_atan_w_lg_w_lg_indexbit10174w10175w(i) <= wire_cata_12_cordic_atan_w_lg_indexbit10174w(0) AND wire_cata_12_cordic_atan_w_valuenode_12_w_range10173w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_12_cordic_atan_w_lg_indexbit10172w(i) <= indexbit AND wire_cata_12_cordic_atan_w_valuenode_15_w_range10171w(i);
	END GENERATE loop7;
	wire_cata_12_cordic_atan_w_lg_indexbit10174w(0) <= NOT indexbit;
	arctan <= (wire_cata_12_cordic_atan_w_lg_w_lg_indexbit10174w10175w OR wire_cata_12_cordic_atan_w_lg_indexbit10172w);
	valuenode_12_w <= "000000000000001111111111111111111111111010101011";
	valuenode_15_w <= "000000000000000001111111111111111111111111111111";
	wire_cata_12_cordic_atan_w_valuenode_12_w_range10173w <= valuenode_12_w(47 DOWNTO 16);
	wire_cata_12_cordic_atan_w_valuenode_15_w_range10171w <= valuenode_15_w(44 DOWNTO 13);

 END RTL; --coshw_altfp_sincos_cordic_atan_m6b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=13 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_n6b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_n6b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_n6b IS

	 SIGNAL  wire_cata_13_cordic_atan_w_lg_w_lg_indexbit10180w10181w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_w_lg_indexbit10178w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_w_lg_indexbit10180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_13_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_16_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_w_valuenode_13_w_range10179w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_w_valuenode_16_w_range10177w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop8 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_13_cordic_atan_w_lg_w_lg_indexbit10180w10181w(i) <= wire_cata_13_cordic_atan_w_lg_indexbit10180w(0) AND wire_cata_13_cordic_atan_w_valuenode_13_w_range10179w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_13_cordic_atan_w_lg_indexbit10178w(i) <= indexbit AND wire_cata_13_cordic_atan_w_valuenode_16_w_range10177w(i);
	END GENERATE loop9;
	wire_cata_13_cordic_atan_w_lg_indexbit10180w(0) <= NOT indexbit;
	arctan <= (wire_cata_13_cordic_atan_w_lg_w_lg_indexbit10180w10181w OR wire_cata_13_cordic_atan_w_lg_indexbit10178w);
	valuenode_13_w <= "000000000000000111111111111111111111111111010101";
	valuenode_16_w <= "000000000000000001000000000000000000000000000000";
	wire_cata_13_cordic_atan_w_valuenode_13_w_range10179w <= valuenode_13_w(47 DOWNTO 16);
	wire_cata_13_cordic_atan_w_valuenode_16_w_range10177w <= valuenode_16_w(44 DOWNTO 13);

 END RTL; --coshw_altfp_sincos_cordic_atan_n6b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=1 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_45b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_45b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_45b IS

	 SIGNAL  wire_cata_1_cordic_atan_w_lg_w_lg_indexbit10186w10187w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_w_lg_indexbit10184w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_w_lg_indexbit10186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_1_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_4_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_w_valuenode_1_w_range10185w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_w_valuenode_4_w_range10183w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop10 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_1_cordic_atan_w_lg_w_lg_indexbit10186w10187w(i) <= wire_cata_1_cordic_atan_w_lg_indexbit10186w(0) AND wire_cata_1_cordic_atan_w_valuenode_1_w_range10185w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_1_cordic_atan_w_lg_indexbit10184w(i) <= indexbit AND wire_cata_1_cordic_atan_w_valuenode_4_w_range10183w(i);
	END GENERATE loop11;
	wire_cata_1_cordic_atan_w_lg_indexbit10186w(0) <= NOT indexbit;
	arctan <= (wire_cata_1_cordic_atan_w_lg_w_lg_indexbit10186w10187w OR wire_cata_1_cordic_atan_w_lg_indexbit10184w);
	valuenode_1_w <= "000111011010110001100111000001010110000110111011";
	valuenode_4_w <= "000000111111111010101011011101101110010110100000";
	wire_cata_1_cordic_atan_w_valuenode_1_w_range10185w <= valuenode_1_w(47 DOWNTO 16);
	wire_cata_1_cordic_atan_w_valuenode_4_w_range10183w <= valuenode_4_w(44 DOWNTO 13);

 END RTL; --coshw_altfp_sincos_cordic_atan_45b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=2 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_55b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_55b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_55b IS

	 SIGNAL  wire_cata_2_cordic_atan_w_lg_w_lg_indexbit10192w10193w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_w_lg_indexbit10190w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_w_lg_indexbit10192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_2_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_5_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_w_valuenode_2_w_range10191w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_w_valuenode_5_w_range10189w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop12 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_2_cordic_atan_w_lg_w_lg_indexbit10192w10193w(i) <= wire_cata_2_cordic_atan_w_lg_indexbit10192w(0) AND wire_cata_2_cordic_atan_w_valuenode_2_w_range10191w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_2_cordic_atan_w_lg_indexbit10190w(i) <= indexbit AND wire_cata_2_cordic_atan_w_valuenode_5_w_range10189w(i);
	END GENERATE loop13;
	wire_cata_2_cordic_atan_w_lg_indexbit10192w(0) <= NOT indexbit;
	arctan <= (wire_cata_2_cordic_atan_w_lg_w_lg_indexbit10192w10193w OR wire_cata_2_cordic_atan_w_lg_indexbit10190w);
	valuenode_2_w <= "000011111010110110111010111111001001011001000000";
	valuenode_5_w <= "000000011111111111010101010110111011101010010111";
	wire_cata_2_cordic_atan_w_valuenode_2_w_range10191w <= valuenode_2_w(47 DOWNTO 16);
	wire_cata_2_cordic_atan_w_valuenode_5_w_range10189w <= valuenode_5_w(44 DOWNTO 13);

 END RTL; --coshw_altfp_sincos_cordic_atan_55b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=3 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_65b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_65b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_65b IS

	 SIGNAL  wire_cata_3_cordic_atan_w_lg_w_lg_indexbit10198w10199w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_w_lg_indexbit10196w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_w_lg_indexbit10198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_3_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_6_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_w_valuenode_3_w_range10197w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_w_valuenode_6_w_range10195w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop14 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_3_cordic_atan_w_lg_w_lg_indexbit10198w10199w(i) <= wire_cata_3_cordic_atan_w_lg_indexbit10198w(0) AND wire_cata_3_cordic_atan_w_valuenode_3_w_range10197w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_3_cordic_atan_w_lg_indexbit10196w(i) <= indexbit AND wire_cata_3_cordic_atan_w_valuenode_6_w_range10195w(i);
	END GENERATE loop15;
	wire_cata_3_cordic_atan_w_lg_indexbit10198w(0) <= NOT indexbit;
	arctan <= (wire_cata_3_cordic_atan_w_lg_w_lg_indexbit10198w10199w OR wire_cata_3_cordic_atan_w_lg_indexbit10196w);
	valuenode_3_w <= "000001111111010101101110101001101010101100001100";
	valuenode_6_w <= "000000001111111111111010101010101101110111011100";
	wire_cata_3_cordic_atan_w_valuenode_3_w_range10197w <= valuenode_3_w(47 DOWNTO 16);
	wire_cata_3_cordic_atan_w_valuenode_6_w_range10195w <= valuenode_6_w(44 DOWNTO 13);

 END RTL; --coshw_altfp_sincos_cordic_atan_65b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=4 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_75b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_75b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_75b IS

	 SIGNAL  wire_cata_4_cordic_atan_w_lg_w_lg_indexbit10204w10205w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_w_lg_indexbit10202w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_w_lg_indexbit10204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_4_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_7_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_w_valuenode_4_w_range10203w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_w_valuenode_7_w_range10201w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop16 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_4_cordic_atan_w_lg_w_lg_indexbit10204w10205w(i) <= wire_cata_4_cordic_atan_w_lg_indexbit10204w(0) AND wire_cata_4_cordic_atan_w_valuenode_4_w_range10203w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_4_cordic_atan_w_lg_indexbit10202w(i) <= indexbit AND wire_cata_4_cordic_atan_w_valuenode_7_w_range10201w(i);
	END GENERATE loop17;
	wire_cata_4_cordic_atan_w_lg_indexbit10204w(0) <= NOT indexbit;
	arctan <= (wire_cata_4_cordic_atan_w_lg_w_lg_indexbit10204w10205w OR wire_cata_4_cordic_atan_w_lg_indexbit10202w);
	valuenode_4_w <= "000000111111111010101011011101101110010110100000";
	valuenode_7_w <= "000000000111111111111111010101010101011011101111";
	wire_cata_4_cordic_atan_w_valuenode_4_w_range10203w <= valuenode_4_w(47 DOWNTO 16);
	wire_cata_4_cordic_atan_w_valuenode_7_w_range10201w <= valuenode_7_w(44 DOWNTO 13);

 END RTL; --coshw_altfp_sincos_cordic_atan_75b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=5 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_85b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_85b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_85b IS

	 SIGNAL  wire_cata_5_cordic_atan_w_lg_w_lg_indexbit10210w10211w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_w_lg_indexbit10208w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_w_lg_indexbit10210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_5_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_8_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_w_valuenode_5_w_range10209w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_w_valuenode_8_w_range10207w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop18 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_5_cordic_atan_w_lg_w_lg_indexbit10210w10211w(i) <= wire_cata_5_cordic_atan_w_lg_indexbit10210w(0) AND wire_cata_5_cordic_atan_w_valuenode_5_w_range10209w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_5_cordic_atan_w_lg_indexbit10208w(i) <= indexbit AND wire_cata_5_cordic_atan_w_valuenode_8_w_range10207w(i);
	END GENERATE loop19;
	wire_cata_5_cordic_atan_w_lg_indexbit10210w(0) <= NOT indexbit;
	arctan <= (wire_cata_5_cordic_atan_w_lg_w_lg_indexbit10210w10211w OR wire_cata_5_cordic_atan_w_lg_indexbit10208w);
	valuenode_5_w <= "000000011111111111010101010110111011101010010111";
	valuenode_8_w <= "000000000011111111111111111010101010101010110111";
	wire_cata_5_cordic_atan_w_valuenode_5_w_range10209w <= valuenode_5_w(47 DOWNTO 16);
	wire_cata_5_cordic_atan_w_valuenode_8_w_range10207w <= valuenode_8_w(44 DOWNTO 13);

 END RTL; --coshw_altfp_sincos_cordic_atan_85b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=6 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_95b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_95b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_95b IS

	 SIGNAL  wire_cata_6_cordic_atan_w_lg_w_lg_indexbit10216w10217w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_w_lg_indexbit10214w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_w_lg_indexbit10216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_6_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_9_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_w_valuenode_6_w_range10215w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_w_valuenode_9_w_range10213w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop20 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_6_cordic_atan_w_lg_w_lg_indexbit10216w10217w(i) <= wire_cata_6_cordic_atan_w_lg_indexbit10216w(0) AND wire_cata_6_cordic_atan_w_valuenode_6_w_range10215w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_6_cordic_atan_w_lg_indexbit10214w(i) <= indexbit AND wire_cata_6_cordic_atan_w_valuenode_9_w_range10213w(i);
	END GENERATE loop21;
	wire_cata_6_cordic_atan_w_lg_indexbit10216w(0) <= NOT indexbit;
	arctan <= (wire_cata_6_cordic_atan_w_lg_w_lg_indexbit10216w10217w OR wire_cata_6_cordic_atan_w_lg_indexbit10214w);
	valuenode_6_w <= "000000001111111111111010101010101101110111011100";
	valuenode_9_w <= "000000000001111111111111111111010101010101010110";
	wire_cata_6_cordic_atan_w_valuenode_6_w_range10215w <= valuenode_6_w(47 DOWNTO 16);
	wire_cata_6_cordic_atan_w_valuenode_9_w_range10213w <= valuenode_9_w(44 DOWNTO 13);

 END RTL; --coshw_altfp_sincos_cordic_atan_95b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=7 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_a5b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_a5b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_a5b IS

	 SIGNAL  wire_cata_7_cordic_atan_w_lg_w_lg_indexbit10222w10223w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_w_lg_indexbit10220w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_w_lg_indexbit10222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_10_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_7_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_w_valuenode_10_w_range10219w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_w_valuenode_7_w_range10221w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop22 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_7_cordic_atan_w_lg_w_lg_indexbit10222w10223w(i) <= wire_cata_7_cordic_atan_w_lg_indexbit10222w(0) AND wire_cata_7_cordic_atan_w_valuenode_7_w_range10221w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_7_cordic_atan_w_lg_indexbit10220w(i) <= indexbit AND wire_cata_7_cordic_atan_w_valuenode_10_w_range10219w(i);
	END GENERATE loop23;
	wire_cata_7_cordic_atan_w_lg_indexbit10222w(0) <= NOT indexbit;
	arctan <= (wire_cata_7_cordic_atan_w_lg_w_lg_indexbit10222w10223w OR wire_cata_7_cordic_atan_w_lg_indexbit10220w);
	valuenode_10_w <= "000000000000111111111111111111111010101010101011";
	valuenode_7_w <= "000000000111111111111111010101010101011011101111";
	wire_cata_7_cordic_atan_w_valuenode_10_w_range10219w <= valuenode_10_w(44 DOWNTO 13);
	wire_cata_7_cordic_atan_w_valuenode_7_w_range10221w <= valuenode_7_w(47 DOWNTO 16);

 END RTL; --coshw_altfp_sincos_cordic_atan_a5b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=8 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_b5b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_b5b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_b5b IS

	 SIGNAL  wire_cata_8_cordic_atan_w_lg_w_lg_indexbit10228w10229w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_w_lg_indexbit10226w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_w_lg_indexbit10228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_11_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_8_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_w_valuenode_11_w_range10225w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_w_valuenode_8_w_range10227w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop24 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_8_cordic_atan_w_lg_w_lg_indexbit10228w10229w(i) <= wire_cata_8_cordic_atan_w_lg_indexbit10228w(0) AND wire_cata_8_cordic_atan_w_valuenode_8_w_range10227w(i);
	END GENERATE loop24;
	loop25 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_8_cordic_atan_w_lg_indexbit10226w(i) <= indexbit AND wire_cata_8_cordic_atan_w_valuenode_11_w_range10225w(i);
	END GENERATE loop25;
	wire_cata_8_cordic_atan_w_lg_indexbit10228w(0) <= NOT indexbit;
	arctan <= (wire_cata_8_cordic_atan_w_lg_w_lg_indexbit10228w10229w OR wire_cata_8_cordic_atan_w_lg_indexbit10226w);
	valuenode_11_w <= "000000000000011111111111111111111111010101010101";
	valuenode_8_w <= "000000000011111111111111111010101010101010110111";
	wire_cata_8_cordic_atan_w_valuenode_11_w_range10225w <= valuenode_11_w(44 DOWNTO 13);
	wire_cata_8_cordic_atan_w_valuenode_8_w_range10227w <= valuenode_8_w(47 DOWNTO 16);

 END RTL; --coshw_altfp_sincos_cordic_atan_b5b


--altfp_sincos_cordic_atan CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" indexpoint=3 START=9 WIDTH=32 arctan indexbit
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_atan_c5b IS 
	 PORT 
	 ( 
		 arctan	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 indexbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_atan_c5b;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_atan_c5b IS

	 SIGNAL  wire_cata_9_cordic_atan_w_lg_w_lg_indexbit10234w10235w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_w_lg_indexbit10232w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_w_lg_indexbit10234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  valuenode_12_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  valuenode_9_w :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_w_valuenode_12_w_range10231w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_w_valuenode_9_w_range10233w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
 BEGIN

	loop26 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_9_cordic_atan_w_lg_w_lg_indexbit10234w10235w(i) <= wire_cata_9_cordic_atan_w_lg_indexbit10234w(0) AND wire_cata_9_cordic_atan_w_valuenode_9_w_range10233w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 31 GENERATE 
		wire_cata_9_cordic_atan_w_lg_indexbit10232w(i) <= indexbit AND wire_cata_9_cordic_atan_w_valuenode_12_w_range10231w(i);
	END GENERATE loop27;
	wire_cata_9_cordic_atan_w_lg_indexbit10234w(0) <= NOT indexbit;
	arctan <= (wire_cata_9_cordic_atan_w_lg_w_lg_indexbit10234w10235w OR wire_cata_9_cordic_atan_w_lg_indexbit10232w);
	valuenode_12_w <= "000000000000001111111111111111111111111010101011";
	valuenode_9_w <= "000000000001111111111111111111010101010101010110";
	wire_cata_9_cordic_atan_w_valuenode_12_w_range10231w <= valuenode_12_w(44 DOWNTO 13);
	wire_cata_9_cordic_atan_w_valuenode_9_w_range10233w <= valuenode_9_w(47 DOWNTO 16);

 END RTL; --coshw_altfp_sincos_cordic_atan_c5b


--altfp_sincos_cordic_start CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" WIDTH=32 index value
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_mux 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_start_509 IS 
	 PORT 
	 ( 
		 index	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
		 value	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END coshw_altfp_sincos_cordic_start_509;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_start_509 IS

	 SIGNAL  wire_mux1_data	:	STD_LOGIC_VECTOR (511 DOWNTO 0);
	 SIGNAL  wire_mux1_data_2d	:	STD_LOGIC_2D(15 DOWNTO 0, 31 DOWNTO 0);
	 SIGNAL  wire_mux1_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  valuenode_0_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_10_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_11_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_12_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_13_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_14_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_15_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_1_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_2_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_3_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_4_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_5_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_6_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_7_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_8_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  valuenode_9_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
 BEGIN

	value <= wire_mux1_result;
	valuenode_0_w <= "001001101101110100111011011010100001";
	valuenode_10_w <= "001111111111111111111101010101010101";
	valuenode_11_w <= "001111111111111111111111010101010101";
	valuenode_12_w <= "001111111111111111111111111101010101";
	valuenode_13_w <= "001111111111111111111111110101010101";
	valuenode_14_w <= "001111111111111111111111111111110101";
	valuenode_15_w <= "001111111111111111111111111111010101";
	valuenode_1_w <= "001101101111011001010110110001011010";
	valuenode_2_w <= "001111010111001100011101111111111011";
	valuenode_3_w <= "001111110101011101000011101100100100";
	valuenode_4_w <= "001111111101010101110100100001100000";
	valuenode_5_w <= "001111111111010101010111010010011001";
	valuenode_6_w <= "001111111111110101010101011101001010";
	valuenode_7_w <= "001111111111111101010101010101110101";
	valuenode_8_w <= "001111111111111111010101010101010111";
	valuenode_9_w <= "001111111111111111110101010101010101";
	wire_mux1_data <= ( valuenode_15_w(35 DOWNTO 4) & valuenode_14_w(35 DOWNTO 4) & valuenode_13_w(35 DOWNTO 4) & valuenode_12_w(35 DOWNTO 4) & valuenode_11_w(35 DOWNTO 4) & valuenode_10_w(35 DOWNTO 4) & valuenode_9_w(35 DOWNTO 4) & valuenode_8_w(35 DOWNTO 4) & valuenode_7_w(35 DOWNTO 4) & valuenode_6_w(35 DOWNTO 4) & valuenode_5_w(35 DOWNTO 4) & valuenode_4_w(35 DOWNTO 4) & valuenode_3_w(35 DOWNTO 4) & valuenode_2_w(35 DOWNTO 4) & valuenode_1_w(35 DOWNTO 4) & valuenode_0_w(35 DOWNTO 4));
	loop28 : FOR i IN 0 TO 15 GENERATE
		loop29 : FOR j IN 0 TO 31 GENERATE
			wire_mux1_data_2d(i, j) <= wire_mux1_data(i*32+j);
		END GENERATE loop29;
	END GENERATE loop28;
	mux1 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 16,
		LPM_WIDTH => 32,
		LPM_WIDTHS => 4
	  )
	  PORT MAP ( 
		data => wire_mux1_data_2d,
		result => wire_mux1_result,
		sel => index
	  );

 END RTL; --coshw_altfp_sincos_cordic_start_509

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 39 lpm_mult 1 lpm_mux 1 reg 1506 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_cordic_m_d5e IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 indexbit	:	IN  STD_LOGIC := '0';
		 radians	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
		 sincos	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 sincosbit	:	IN  STD_LOGIC := '0'
	 ); 
 END coshw_altfp_sincos_cordic_m_d5e;

 ARCHITECTURE RTL OF coshw_altfp_sincos_cordic_m_d5e IS

	 SIGNAL  wire_cata_0_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_10_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_11_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_12_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_13_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_1_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_2_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_3_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_4_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_5_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_6_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_7_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_8_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cata_9_cordic_atan_arctan	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cxs_value	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 cdaff_0	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cdaff_1	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cdaff_2	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 indexbitff	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_indexbitff_w_lg_w_q_range448w546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range477w7967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range480w8718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range483w9464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range9992w9995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range450w983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range453w1779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range456w2570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range459w3356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range462w4137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range465w4913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range468w5684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range471w6450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_lg_w_q_range474w7211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range9992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_indexbitff_w_q_range474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 sincosbitff	:	STD_LOGIC_VECTOR(16 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_sincosbitff_w_lg_w_q_range535w9982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sincosbitff_w_lg_w_q_range9989w9990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sincosbitff_w_q_range535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sincosbitff_w_q_range9989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 sincosff	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_0	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range547w548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range584w601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range584w585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range589w606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range589w590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range594w611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range594w595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range599w616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range599w600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range604w621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range604w605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range609w626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range609w610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range614w631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range614w615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range619w636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range619w620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range624w641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range624w625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range629w646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range629w630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range554w555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range634w651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range634w635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range639w656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range639w640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range644w661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range644w645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range649w666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range649w650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range654w671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range654w655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range659w676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range659w660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range664w681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range664w665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range669w686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range669w670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range674w691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range674w675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range679w694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range679w680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range560w561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range684w696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range684w685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range689w690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range544w566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range544w545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range552w571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range552w553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range558w576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range558w559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range564w581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range564w565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range569w586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range569w570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range574w591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range574w575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range579w596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range579w580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_q_range689w698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range547w548w549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range584w601w602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range589w606w607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range594w611w612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range599w616w617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range604w621w622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range609w626w627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range614w631w632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range619w636w637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range624w641w642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range629w646w647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range554w555w556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range634w651w652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range639w656w657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range644w661w662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range649w666w667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range654w671w672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range659w676w677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range664w681w682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range669w686w687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range674w691w692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range560w561w562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range544w566w567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range552w571w572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range558w576w577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range564w581w582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range569w586w587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range574w591w592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_lg_w_lg_w_q_range579w596w597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_0_w_q_range579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 x_pipeff_1	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_10	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_11	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_12	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_13	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_x_pipeff_13_w_lg_q9987w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_x_pipeff_13_w_lg_q9984w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 x_pipeff_2	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_3	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_4	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_5	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_6	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_7	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_8	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 x_pipeff_9	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 y_pipeff_0	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 y_pipeff_1	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range770w771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range776w777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range782w783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range788w789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range794w795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range800w801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range806w807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range812w813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range818w819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range824w825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range717w718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range830w831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range836w837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range842w843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range848w849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range854w855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range860w861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range866w867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range872w873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range878w879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range884w885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range722w723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range890w891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range700w701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range728w729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range734w735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range740w741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range746w747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range752w753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range758w759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_lg_w_q_range764w765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_1_w_q_range764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_10	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7782w7783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7787w7788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7793w7794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7799w7800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7805w7806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7811w7812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7817w7818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7823w7824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7829w7830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7835w7836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7841w7842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7847w7848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7853w7854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7859w7860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7865w7866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7871w7872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7877w7878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7883w7884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7889w7890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7895w7896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7901w7902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_lg_w_q_range7729w7730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_10_w_q_range7729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_11	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8542w8543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8547w8548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8553w8554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8559w8560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8565w8566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8571w8572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8577w8578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8583w8584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8589w8590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8595w8596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8601w8602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8607w8608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8613w8614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8619w8620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8625w8626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8631w8632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8637w8638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8643w8644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8649w8650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8655w8656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_lg_w_q_range8485w8486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_11_w_q_range8485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_12	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9297w9298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9302w9303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9308w9309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9314w9315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9320w9321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9326w9327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9332w9333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9338w9339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9344w9345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9350w9351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9356w9357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9362w9363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9368w9369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9374w9375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9380w9381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9386w9387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9392w9393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9398w9399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9404w9405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_lg_w_q_range9236w9237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_12_w_q_range9236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_13	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_13_w_lg_q9983w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_13_w_lg_q9986w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 y_pipeff_2	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1569w1570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1575w1576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1581w1582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1587w1588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1593w1594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1599w1600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1605w1606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1611w1612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1617w1618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1623w1624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1629w1630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1635w1636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1641w1642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1647w1648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1653w1654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1659w1660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1665w1666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1671w1672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1677w1678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1683w1684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1522w1523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1689w1690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1501w1502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1527w1528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1533w1534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1539w1540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1545w1546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1551w1552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1557w1558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_lg_w_q_range1563w1564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_2_w_q_range1563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_3	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2363w2364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2369w2370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2375w2376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2381w2382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2387w2388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2393w2394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2399w2400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2405w2406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2411w2412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2417w2418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2423w2424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2429w2430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2435w2436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2441w2442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2447w2448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2453w2454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2459w2460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2465w2466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2471w2472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2477w2478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2483w2484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2297w2298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2322w2323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2327w2328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2333w2334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2339w2340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2345w2346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2351w2352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_lg_w_q_range2357w2358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_3_w_q_range2357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_4	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3152w3153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3158w3159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3164w3165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3170w3171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3176w3177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3182w3183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3188w3189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3194w3195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3200w3201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3206w3207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3212w3213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3218w3219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3224w3225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3230w3231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3236w3237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3242w3243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3248w3249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3254w3255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3260w3261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3266w3267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3272w3273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3088w3089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3117w3118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3122w3123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3128w3129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3134w3135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3140w3141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_lg_w_q_range3146w3147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_4_w_q_range3146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_5	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3936w3937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3942w3943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3948w3949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3954w3955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3960w3961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3966w3967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3972w3973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3978w3979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3984w3985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3990w3991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3996w3997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4002w4003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4008w4009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4014w4015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4020w4021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4026w4027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4032w4033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4038w4039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4044w4045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4050w4051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range4056w4057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3874w3875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3907w3908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3912w3913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3918w3919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3924w3925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_lg_w_q_range3930w3931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range4056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_5_w_q_range3930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_6	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4715w4716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4721w4722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4727w4728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4733w4734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4739w4740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4745w4746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4751w4752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4757w4758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4763w4764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4769w4770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4775w4776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4781w4782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4787w4788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4793w4794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4799w4800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4805w4806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4811w4812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4817w4818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4823w4824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4829w4830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4835w4836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4655w4656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4692w4693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4697w4698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4703w4704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_lg_w_q_range4709w4710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_6_w_q_range4709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_7	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5489w5490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5495w5496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5501w5502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5507w5508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5513w5514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5519w5520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5525w5526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5531w5532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5537w5538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5543w5544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5549w5550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5555w5556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5561w5562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5567w5568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5573w5574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5579w5580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5585w5586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5591w5592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5597w5598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5603w5604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5609w5610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5431w5432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5472w5473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5477w5478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_lg_w_q_range5483w5484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_7_w_q_range5483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_8	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6258w6259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6264w6265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6270w6271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6276w6277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6282w6283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6288w6289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6294w6295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6300w6301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6306w6307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6312w6313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6318w6319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6324w6325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6330w6331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6336w6337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6342w6343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6348w6349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6354w6355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6360w6361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6366w6367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6372w6373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6378w6379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6202w6203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6247w6248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_lg_w_q_range6252w6253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_8_w_q_range6252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 y_pipeff_9	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7022w7023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7028w7029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7034w7035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7040w7041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7046w7047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7052w7053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7058w7059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7064w7065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7070w7071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7076w7077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7082w7083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7088w7089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7094w7095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7100w7101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7106w7107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7112w7113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7118w7119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7124w7125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7130w7131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7136w7137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7142w7143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range6968w6969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_lg_w_q_range7017w7018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range6968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_y_pipeff_9_w_q_range7017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_0	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 z_pipeff_1	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_1_w_q_range1241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_10	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_10_w_q_range8225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_11	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_11_w_q_range8976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_12	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_12_w_q_range9722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_13	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 z_pipeff_2	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_2_w_q_range2037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_3	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_3_w_q_range2828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_4	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_4_w_q_range3614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_5	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_5_w_q_range4395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_6	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_6_w_q_range5171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_7	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_7_w_q_range5942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_8	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_8_w_q_range6708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 z_pipeff_9	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_z_pipeff_9_w_q_range7469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_sincos_add_cin	:	STD_LOGIC;
	 SIGNAL  wire_sincos_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_10_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_11_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_12_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_13_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_2_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_3_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_4_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_5_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_6_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_7_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_8_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_x_pipenode_9_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipeff1_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_10_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_11_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_12_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_13_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_2_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_3_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_4_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_5_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_6_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_7_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_8_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_y_pipenode_9_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_z_pipeff1_sub_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_10_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_11_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_12_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_13_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_2_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_3_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_4_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_5_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_6_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_7_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_8_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_z_pipenode_9_add_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_cmx_result	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_indexpointnum_w288w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range9996w9997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10033w10050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10033w10034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10038w10055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10038w10039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10043w10060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10043w10044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10048w10065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10048w10049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10053w10070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10053w10054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10058w10075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10058w10059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10063w10080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10063w10064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10068w10085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10068w10069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10073w10090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10073w10074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10078w10095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10078w10079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10003w10004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10083w10100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10083w10084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10088w10105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10088w10089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10093w10110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10093w10094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10098w10115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10098w10099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10103w10120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10103w10104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10108w10125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10108w10109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10113w10130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10113w10114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10118w10135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10118w10119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10123w10140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10123w10124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10128w10143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10128w10129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10009w10010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10133w10146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10133w10134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10138w10149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10138w10139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range9993w10015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range9993w9994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10001w10020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10001w10002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10007w10025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10007w10008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10013w10030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10013w10014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10018w10035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10018w10019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10023w10040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10023w10024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10028w10045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10028w10029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range289w292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range289w302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range335w338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range335w352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range340w343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range340w357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range345w348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range345w362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range350w353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range350w367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range355w358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range355w372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range360w363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range360w377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range365w368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range365w382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range370w373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range370w387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range375w378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range375w392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range380w383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range380w397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range294w296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range294w307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range385w388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range385w402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range390w393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range390w407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range395w398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range395w412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range400w403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range400w417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range405w408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range405w422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range410w413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range410w427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range415w418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range415w432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range420w423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range420w437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range425w428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range425w442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range430w433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range297w299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range297w312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range435w438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range440w443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range300w303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range300w317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range305w308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range305w322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range310w313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range310w327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range315w318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range315w332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range320w323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range320w337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range325w328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range325w342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range330w333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_radians_range330w347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7019w7212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7078w7294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7084w7302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7090w7310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7096w7318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7102w7326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7108w7334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7114w7342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7120w7350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7126w7358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7132w7366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7024w7222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7138w7374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7144w7382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7148w7390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6970w7398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6975w7406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6977w7414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6979w7422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6981w7430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6983w7438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6985w7446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7030w7230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6987w7454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6989w7462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7036w7238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7042w7246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7048w7254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7054w7262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7060w7270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7066w7278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7072w7286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7784w7968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7843w8050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7849w8058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7855w8066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7861w8074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7867w8082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7873w8090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7879w8098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7885w8106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7891w8114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7897w8122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7789w7978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7903w8130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7907w8138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7731w8146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7736w8154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7738w8162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7740w8170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7742w8178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7744w8186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7746w8194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7748w8202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7795w7986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7750w8210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7752w8218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7801w7994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7807w8002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7813w8010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7819w8018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7825w8026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7831w8034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7837w8042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8544w8719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8603w8801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8609w8809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8615w8817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8621w8825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8627w8833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8633w8841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8639w8849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8645w8857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8651w8865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8657w8873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8549w8729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8661w8881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8487w8889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8492w8897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8494w8905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8496w8913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8498w8921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8500w8929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8502w8937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8504w8945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8506w8953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8555w8737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8508w8961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8510w8969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8561w8745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8567w8753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8573w8761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8579w8769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8585w8777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8591w8785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8597w8793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9299w9465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9358w9547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9364w9555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9370w9563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9376w9571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9382w9579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9388w9587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9394w9595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9400w9603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9406w9611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9410w9619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9304w9475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9238w9627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9243w9635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9245w9643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9247w9651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9249w9659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9251w9667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9253w9675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9255w9683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9257w9691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9259w9699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9310w9483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9261w9707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9263w9715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9316w9491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9322w9499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9328w9507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9334w9515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9340w9523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9346w9531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9352w9539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range719w984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range778w1066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range784w1074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range790w1082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range796w1090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range802w1098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range808w1106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range814w1114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range820w1122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range826w1130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range832w1138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range724w994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range838w1146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range844w1154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range850w1162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range856w1170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range862w1178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range868w1186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range874w1194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range880w1202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range886w1210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range892w1218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range730w1002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range896w1226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range702w1234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range736w1010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range742w1018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range748w1026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range754w1034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range760w1042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range766w1050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range772w1058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1524w1780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1583w1862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1589w1870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1595w1878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1601w1886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1607w1894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1613w1902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1619w1910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1625w1918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1631w1926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1637w1934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1529w1790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1643w1942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1649w1950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1655w1958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1661w1966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1667w1974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1673w1982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1679w1990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1685w1998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1691w2006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1695w2014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1535w1798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1503w2022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1508w2030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1541w1806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1547w1814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1553w1822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1559w1830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1565w1838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1571w1846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1577w1854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2324w2571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2383w2653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2389w2661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2395w2669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2401w2677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2407w2685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2413w2693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2419w2701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2425w2709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2431w2717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2437w2725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2329w2581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2443w2733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2449w2741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2455w2749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2461w2757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2467w2765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2473w2773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2479w2781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2485w2789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2489w2797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2299w2805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2335w2589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2304w2813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2306w2821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2341w2597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2347w2605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2353w2613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2359w2621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2365w2629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2371w2637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2377w2645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3119w3357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3178w3439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3184w3447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3190w3455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3196w3463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3202w3471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3208w3479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3214w3487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3220w3495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3226w3503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3232w3511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3124w3367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3238w3519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3244w3527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3250w3535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3256w3543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3262w3551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3268w3559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3274w3567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3278w3575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3090w3583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3095w3591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3130w3375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3097w3599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3099w3607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3136w3383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3142w3391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3148w3399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3154w3407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3160w3415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3166w3423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3172w3431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3909w4138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3968w4220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3974w4228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3980w4236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3986w4244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3992w4252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3998w4260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4004w4268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4010w4276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4016w4284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4022w4292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3914w4148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4028w4300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4034w4308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4040w4316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4046w4324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4052w4332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4058w4340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4062w4348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3876w4356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3881w4364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3883w4372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3920w4156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3885w4380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3887w4388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3926w4164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3932w4172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3938w4180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3944w4188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3950w4196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3956w4204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3962w4212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4694w4914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4753w4996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4759w5004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4765w5012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4771w5020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4777w5028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4783w5036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4789w5044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4795w5052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4801w5060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4807w5068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4699w4924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4813w5076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4819w5084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4825w5092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4831w5100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4837w5108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4841w5116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4657w5124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4662w5132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4664w5140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4666w5148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4705w4932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4668w5156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4670w5164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4711w4940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4717w4948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4723w4956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4729w4964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4735w4972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4741w4980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4747w4988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5474w5685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5533w5767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5539w5775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5545w5783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5551w5791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5557w5799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5563w5807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5569w5815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5575w5823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5581w5831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5587w5839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5479w5695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5593w5847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5599w5855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5605w5863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5611w5871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5615w5879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5433w5887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5438w5895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5440w5903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5442w5911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5444w5919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5485w5703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5446w5927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5448w5935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5491w5711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5497w5719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5503w5727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5509w5735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5515w5743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5521w5751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5527w5759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6249w6451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6308w6533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6314w6541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6320w6549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6326w6557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6332w6565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6338w6573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6344w6581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6350w6589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6356w6597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6362w6605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6254w6461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6368w6613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6374w6621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6380w6629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6384w6637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6204w6645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6209w6653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6211w6661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6213w6669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6215w6677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6217w6685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6260w6469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6219w6693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6221w6701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6266w6477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6272w6485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6278w6493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6284w6501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6290w6509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6296w6517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6302w6525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7151w7210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7180w7293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7183w7301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7186w7309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7189w7317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7192w7325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7195w7333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7198w7341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7201w7349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7204w7357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7207w7365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7153w7221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range6991w7373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range6995w7381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range6997w7389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range6999w7397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7001w7405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7003w7413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7005w7421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7007w7429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7009w7437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7011w7445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7156w7229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7013w7453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7015w7461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7159w7237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7162w7245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7165w7253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7168w7261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7171w7269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7174w7277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7177w7285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7910w7966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7939w8049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7942w8057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7945w8065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7948w8073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7951w8081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7954w8089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7957w8097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7960w8105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7963w8113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7754w8121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7912w7977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7758w8129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7760w8137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7762w8145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7764w8153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7766w8161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7768w8169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7770w8177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7772w8185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7774w8193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7776w8201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7915w7985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7778w8209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7780w8217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7918w7993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7921w8001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7924w8009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7927w8017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7930w8025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7933w8033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7936w8041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8664w8717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8693w8800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8696w8808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8699w8816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8702w8824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8705w8832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8708w8840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8711w8848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8714w8856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8512w8864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8516w8872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8666w8728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8518w8880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8520w8888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8522w8896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8524w8904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8526w8912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8528w8920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8530w8928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8532w8936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8534w8944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8536w8952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8669w8736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8538w8960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8540w8968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8672w8744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8675w8752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8678w8760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8681w8768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8684w8776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8687w8784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8690w8792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9413w9463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9442w9546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9445w9554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9448w9562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9451w9570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9454w9578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9457w9586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9460w9594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9265w9602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9269w9610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9271w9618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9415w9474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9273w9626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9275w9634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9277w9642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9279w9650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9281w9658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9283w9666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9285w9674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9287w9682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9289w9690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9291w9698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9418w9482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9293w9706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9295w9714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9421w9490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9424w9498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9427w9506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9430w9514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9433w9522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9436w9530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9439w9538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range899w982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range928w1065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range931w1073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range934w1081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range937w1089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range940w1097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range943w1105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range946w1113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range949w1121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range952w1129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range955w1137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range901w993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range958w1145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range961w1153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range964w1161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range967w1169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range970w1177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range973w1185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range976w1193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range979w1201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range707w1209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range711w1217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range904w1001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range713w1225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range715w1233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range907w1009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range910w1017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range913w1025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range916w1033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range919w1041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range922w1049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range925w1057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1698w1778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1727w1861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1730w1869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1733w1877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1736w1885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1739w1893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1742w1901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1745w1909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1748w1917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1751w1925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1754w1933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1700w1789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1757w1941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1760w1949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1763w1957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1766w1965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1769w1973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1772w1981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1775w1989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1510w1997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1514w2005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1516w2013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1703w1797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1518w2021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1520w2029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1706w1805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1709w1813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1712w1821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1715w1829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1718w1837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1721w1845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1724w1853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2492w2569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2521w2652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2524w2660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2527w2668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2530w2676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2533w2684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2536w2692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2539w2700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2542w2708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2545w2716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2548w2724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2494w2580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2551w2732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2554w2740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2557w2748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2560w2756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2563w2764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2566w2772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2308w2780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2312w2788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2314w2796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2316w2804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2497w2588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2318w2812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2320w2820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2500w2596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2503w2604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2506w2612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2509w2620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2512w2628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2515w2636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2518w2644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3281w3355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3310w3438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3313w3446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3316w3454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3319w3462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3322w3470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3325w3478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3328w3486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3331w3494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3334w3502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3337w3510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3283w3366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3340w3518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3343w3526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3346w3534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3349w3542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3352w3550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3101w3558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3105w3566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3107w3574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3109w3582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3111w3590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3286w3374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3113w3598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3115w3606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3289w3382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3292w3390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3295w3398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3298w3406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3301w3414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3304w3422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3307w3430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4065w4136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4094w4219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4097w4227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4100w4235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4103w4243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4106w4251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4109w4259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4112w4267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4115w4275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4118w4283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4121w4291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4067w4147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4124w4299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4127w4307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4130w4315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4133w4323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3889w4331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3893w4339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3895w4347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3897w4355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3899w4363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3901w4371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4070w4155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3903w4379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3905w4387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4073w4163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4076w4171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4079w4179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4082w4187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4085w4195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4088w4203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4091w4211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4844w4912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4873w4995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4876w5003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4879w5011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4882w5019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4885w5027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4888w5035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4891w5043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4894w5051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4897w5059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4900w5067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4846w4923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4903w5075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4906w5083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4909w5091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4672w5099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4676w5107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4678w5115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4680w5123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4682w5131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4684w5139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4686w5147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4849w4931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4688w5155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4690w5163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4852w4939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4855w4947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4858w4955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4861w4963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4864w4971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4867w4979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4870w4987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5618w5683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5647w5766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5650w5774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5653w5782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5656w5790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5659w5798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5662w5806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5665w5814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5668w5822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5671w5830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5674w5838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5620w5694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5677w5846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5680w5854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5450w5862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5454w5870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5456w5878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5458w5886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5460w5894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5462w5902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5464w5910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5466w5918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5623w5702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5468w5926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5470w5934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5626w5710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5629w5718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5632w5726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5635w5734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5638w5742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5641w5750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5644w5758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6387w6449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6416w6532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6419w6540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6422w6548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6425w6556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6428w6564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6431w6572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6434w6580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6437w6588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6440w6596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6443w6604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6389w6460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6446w6612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6223w6620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6227w6628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6229w6636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6231w6644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6233w6652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6235w6660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6237w6668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6239w6676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6241w6684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6392w6468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6243w6692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6245w6700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6395w6476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6398w6484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6401w6492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6404w6500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6407w6508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6410w6516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6413w6524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7021w7217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7080w7298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7086w7306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7092w7314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7098w7322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7104w7330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7110w7338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7116w7346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7122w7354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7128w7362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7134w7370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7026w7226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7140w7378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7146w7386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7149w7394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6973w7402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6976w7410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6978w7418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6980w7426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6982w7434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6984w7442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6986w7450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7032w7234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6988w7458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6990w7466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7038w7242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7044w7250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7050w7258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7056w7266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7062w7274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7068w7282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7074w7290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7786w7973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7845w8054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7851w8062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7857w8070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7863w8078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7869w8086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7875w8094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7881w8102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7887w8110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7893w8118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7899w8126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7791w7982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7905w8134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7908w8142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7734w8150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7737w8158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7739w8166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7741w8174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7743w8182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7745w8190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7747w8198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7749w8206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7797w7990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7751w8214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7753w8222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7803w7998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7809w8006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7815w8014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7821w8022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7827w8030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7833w8038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7839w8046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8546w8724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8605w8805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8611w8813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8617w8821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8623w8829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8629w8837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8635w8845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8641w8853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8647w8861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8653w8869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8659w8877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8551w8733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8662w8885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8490w8893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8493w8901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8495w8909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8497w8917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8499w8925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8501w8933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8503w8941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8505w8949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8507w8957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8557w8741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8509w8965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8511w8973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8563w8749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8569w8757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8575w8765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8581w8773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8587w8781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8593w8789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8599w8797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9301w9470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9360w9551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9366w9559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9372w9567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9378w9575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9384w9583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9390w9591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9396w9599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9402w9607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9408w9615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9411w9623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9306w9479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9241w9631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9244w9639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9246w9647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9248w9655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9250w9663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9252w9671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9254w9679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9256w9687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9258w9695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9260w9703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9312w9487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9262w9711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9264w9719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9318w9495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9324w9503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9330w9511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9336w9519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9342w9527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9348w9535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9354w9543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range721w989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range780w1070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range786w1078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range792w1086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range798w1094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range804w1102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range810w1110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range816w1118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range822w1126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range828w1134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range834w1142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range726w998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range840w1150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range846w1158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range852w1166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range858w1174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range864w1182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range870w1190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range876w1198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range882w1206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range888w1214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range894w1222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range732w1006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range897w1230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range705w1238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range738w1014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range744w1022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range750w1030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range756w1038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range762w1046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range768w1054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range774w1062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1526w1785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1585w1866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1591w1874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1597w1882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1603w1890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1609w1898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1615w1906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1621w1914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1627w1922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1633w1930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1639w1938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1531w1794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1645w1946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1651w1954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1657w1962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1663w1970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1669w1978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1675w1986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1681w1994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1687w2002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1693w2010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1696w2018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1537w1802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1506w2026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1509w2034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1543w1810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1549w1818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1555w1826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1561w1834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1567w1842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1573w1850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1579w1858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2326w2576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2385w2657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2391w2665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2397w2673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2403w2681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2409w2689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2415w2697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2421w2705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2427w2713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2433w2721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2439w2729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2331w2585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2445w2737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2451w2745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2457w2753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2463w2761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2469w2769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2475w2777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2481w2785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2487w2793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2490w2801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2302w2809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2337w2593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2305w2817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2307w2825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2343w2601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2349w2609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2355w2617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2361w2625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2367w2633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2373w2641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2379w2649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3121w3362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3180w3443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3186w3451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3192w3459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3198w3467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3204w3475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3210w3483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3216w3491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3222w3499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3228w3507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3234w3515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3126w3371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3240w3523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3246w3531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3252w3539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3258w3547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3264w3555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3270w3563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3276w3571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3279w3579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3093w3587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3096w3595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3132w3379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3098w3603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3100w3611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3138w3387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3144w3395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3150w3403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3156w3411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3162w3419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3168w3427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3174w3435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3911w4143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3970w4224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3976w4232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3982w4240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3988w4248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3994w4256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4000w4264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4006w4272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4012w4280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4018w4288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4024w4296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3916w4152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4030w4304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4036w4312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4042w4320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4048w4328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4054w4336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4060w4344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4063w4352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3879w4360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3882w4368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3884w4376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3922w4160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3886w4384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3888w4392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3928w4168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3934w4176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3940w4184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3946w4192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3952w4200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3958w4208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3964w4216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4696w4919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4755w5000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4761w5008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4767w5016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4773w5024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4779w5032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4785w5040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4791w5048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4797w5056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4803w5064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4809w5072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4701w4928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4815w5080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4821w5088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4827w5096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4833w5104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4839w5112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4842w5120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4660w5128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4663w5136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4665w5144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4667w5152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4707w4936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4669w5160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4671w5168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4713w4944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4719w4952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4725w4960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4731w4968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4737w4976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4743w4984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4749w4992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5476w5690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5535w5771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5541w5779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5547w5787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5553w5795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5559w5803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5565w5811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5571w5819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5577w5827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5583w5835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5589w5843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5481w5699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5595w5851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5601w5859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5607w5867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5613w5875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5616w5883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5436w5891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5439w5899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5441w5907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5443w5915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5445w5923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5487w5707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5447w5931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5449w5939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5493w5715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5499w5723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5505w5731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5511w5739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5517w5747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5523w5755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5529w5763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6251w6456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6310w6537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6316w6545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6322w6553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6328w6561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6334w6569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6340w6577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6346w6585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6352w6593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6358w6601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6364w6609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6256w6465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6370w6617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6376w6625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6382w6633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6385w6641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6207w6649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6210w6657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6212w6665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6214w6673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6216w6681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6218w6689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6262w6473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6220w6697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6222w6705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6268w6481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6274w6489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6280w6497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6286w6505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6292w6513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6298w6521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6304w6529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7152w7216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7181w7297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7184w7305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7187w7313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7190w7321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7193w7329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7196w7337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7199w7345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7202w7353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7205w7361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7208w7369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7154w7225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range6993w7377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range6996w7385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range6998w7393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7000w7401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7002w7409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7004w7417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7006w7425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7008w7433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7010w7441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7012w7449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7157w7233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7014w7457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7016w7465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7160w7241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7163w7249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7166w7257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7169w7265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7172w7273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7175w7281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7178w7289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7911w7972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7940w8053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7943w8061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7946w8069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7949w8077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7952w8085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7955w8093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7958w8101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7961w8109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7964w8117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7756w8125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7913w7981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7759w8133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7761w8141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7763w8149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7765w8157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7767w8165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7769w8173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7771w8181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7773w8189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7775w8197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7777w8205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7916w7989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7779w8213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7781w8221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7919w7997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7922w8005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7925w8013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7928w8021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7931w8029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7934w8037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7937w8045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8665w8723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8694w8804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8697w8812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8700w8820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8703w8828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8706w8836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8709w8844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8712w8852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8715w8860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8514w8868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8517w8876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8667w8732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8519w8884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8521w8892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8523w8900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8525w8908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8527w8916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8529w8924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8531w8932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8533w8940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8535w8948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8537w8956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8670w8740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8539w8964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8541w8972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8673w8748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8676w8756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8679w8764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8682w8772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8685w8780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8688w8788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8691w8796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9414w9469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9443w9550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9446w9558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9449w9566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9452w9574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9455w9582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9458w9590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9461w9598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9267w9606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9270w9614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9272w9622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9416w9478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9274w9630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9276w9638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9278w9646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9280w9654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9282w9662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9284w9670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9286w9678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9288w9686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9290w9694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9292w9702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9419w9486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9294w9710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9296w9718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9422w9494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9425w9502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9428w9510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9431w9518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9434w9526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9437w9534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9440w9542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range900w988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range929w1069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range932w1077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range935w1085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range938w1093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range941w1101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range944w1109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range947w1117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range950w1125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range953w1133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range956w1141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range902w997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range959w1149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range962w1157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range965w1165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range968w1173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range971w1181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range974w1189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range977w1197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range980w1205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range709w1213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range712w1221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range905w1005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range714w1229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range716w1237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range908w1013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range911w1021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range914w1029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range917w1037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range920w1045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range923w1053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range926w1061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1699w1784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1728w1865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1731w1873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1734w1881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1737w1889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1740w1897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1743w1905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1746w1913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1749w1921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1752w1929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1755w1937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1701w1793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1758w1945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1761w1953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1764w1961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1767w1969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1770w1977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1773w1985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1776w1993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1512w2001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1515w2009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1517w2017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1704w1801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1519w2025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1521w2033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1707w1809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1710w1817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1713w1825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1716w1833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1719w1841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1722w1849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1725w1857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2493w2575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2522w2656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2525w2664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2528w2672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2531w2680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2534w2688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2537w2696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2540w2704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2543w2712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2546w2720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2549w2728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2495w2584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2552w2736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2555w2744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2558w2752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2561w2760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2564w2768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2567w2776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2310w2784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2313w2792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2315w2800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2317w2808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2498w2592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2319w2816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2321w2824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2501w2600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2504w2608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2507w2616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2510w2624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2513w2632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2516w2640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2519w2648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3282w3361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3311w3442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3314w3450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3317w3458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3320w3466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3323w3474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3326w3482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3329w3490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3332w3498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3335w3506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3338w3514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3284w3370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3341w3522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3344w3530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3347w3538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3350w3546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3353w3554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3103w3562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3106w3570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3108w3578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3110w3586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3112w3594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3287w3378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3114w3602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3116w3610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3290w3386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3293w3394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3296w3402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3299w3410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3302w3418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3305w3426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3308w3434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4066w4142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4095w4223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4098w4231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4101w4239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4104w4247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4107w4255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4110w4263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4113w4271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4116w4279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4119w4287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4122w4295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4068w4151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4125w4303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4128w4311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4131w4319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4134w4327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3891w4335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3894w4343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3896w4351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3898w4359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3900w4367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3902w4375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4071w4159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3904w4383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3906w4391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4074w4167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4077w4175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4080w4183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4083w4191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4086w4199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4089w4207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4092w4215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4845w4918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4874w4999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4877w5007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4880w5015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4883w5023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4886w5031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4889w5039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4892w5047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4895w5055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4898w5063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4901w5071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4847w4927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4904w5079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4907w5087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4910w5095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4674w5103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4677w5111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4679w5119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4681w5127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4683w5135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4685w5143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4687w5151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4850w4935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4689w5159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4691w5167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4853w4943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4856w4951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4859w4959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4862w4967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4865w4975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4868w4983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4871w4991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5619w5689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5648w5770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5651w5778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5654w5786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5657w5794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5660w5802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5663w5810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5666w5818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5669w5826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5672w5834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5675w5842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5621w5698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5678w5850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5681w5858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5452w5866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5455w5874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5457w5882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5459w5890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5461w5898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5463w5906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5465w5914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5467w5922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5624w5706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5469w5930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5471w5938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5627w5714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5630w5722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5633w5730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5636w5738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5639w5746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5642w5754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5645w5762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6388w6455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6417w6536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6420w6544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6423w6552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6426w6560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6429w6568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6432w6576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6435w6584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6438w6592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6441w6600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6444w6608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6390w6464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6447w6616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6225w6624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6228w6632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6230w6640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6232w6648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6234w6656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6236w6664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6238w6672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6240w6680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6242w6688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6393w6472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6244w6696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6246w6704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6396w6480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6399w6488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6402w6496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6405w6504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6408w6512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6411w6520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6414w6528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_indexbit291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8232w8233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8313w8314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8321w8322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8329w8330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8337w8338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8345w8346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8353w8354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8361w8362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8369w8370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8377w8378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8385w8386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8241w8242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8393w8394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8401w8402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8409w8410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8417w8418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8425w8426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8433w8434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8441w8442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8449w8450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8457w8458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8465w8466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8249w8250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8473w8474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8481w8482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8257w8258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8265w8266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8273w8274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8281w8282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8289w8290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8297w8298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8305w8306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range8983w8984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9064w9065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9072w9073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9080w9081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9088w9089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9096w9097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9104w9105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9112w9113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9120w9121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9128w9129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9136w9137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range8992w8993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9144w9145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9152w9153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9160w9161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9168w9169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9176w9177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9184w9185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9192w9193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9200w9201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9208w9209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9216w9217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9000w9001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9224w9225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9232w9233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9008w9009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9016w9017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9024w9025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9032w9033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9040w9041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9048w9049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9056w9057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9729w9730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9810w9811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9818w9819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9826w9827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9834w9835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9842w9843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9850w9851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9858w9859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9866w9867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9874w9875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9882w9883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9738w9739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9890w9891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9898w9899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9906w9907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9914w9915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9922w9923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9930w9931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9938w9939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9946w9947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9954w9955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9962w9963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9746w9747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9970w9971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9978w9979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9754w9755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9762w9763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9770w9771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9778w9779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9786w9787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9794w9795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9802w9803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1248w1249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1329w1330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1337w1338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1345w1346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1353w1354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1361w1362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1369w1370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1377w1378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1385w1386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1393w1394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1401w1402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1257w1258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1409w1410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1417w1418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1425w1426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1433w1434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1441w1442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1449w1450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1457w1458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1465w1466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1473w1474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1481w1482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1265w1266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1489w1490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1497w1498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1273w1274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1281w1282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1289w1290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1297w1298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1305w1306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1313w1314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1321w1322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2044w2045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2125w2126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2133w2134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2141w2142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2149w2150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2157w2158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2165w2166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2173w2174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2181w2182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2189w2190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2197w2198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2053w2054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2205w2206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2213w2214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2221w2222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2229w2230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2237w2238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2245w2246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2253w2254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2261w2262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2269w2270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2277w2278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2061w2062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2285w2286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2293w2294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2069w2070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2077w2078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2085w2086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2093w2094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2101w2102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2109w2110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2117w2118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2835w2836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2916w2917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2924w2925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2932w2933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2940w2941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2948w2949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2956w2957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2964w2965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2972w2973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2980w2981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2988w2989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2844w2845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2996w2997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3004w3005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3012w3013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3020w3021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3028w3029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3036w3037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3044w3045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3052w3053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3060w3061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3068w3069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2852w2853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3076w3077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3084w3085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2860w2861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2868w2869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2876w2877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2884w2885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2892w2893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2900w2901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2908w2909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3621w3622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3702w3703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3710w3711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3718w3719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3726w3727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3734w3735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3742w3743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3750w3751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3758w3759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3766w3767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3774w3775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3630w3631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3782w3783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3790w3791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3798w3799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3806w3807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3814w3815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3822w3823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3830w3831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3838w3839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3846w3847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3854w3855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3638w3639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3862w3863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3870w3871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3646w3647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3654w3655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3662w3663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3670w3671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3678w3679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3686w3687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3694w3695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4402w4403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4483w4484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4491w4492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4499w4500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4507w4508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4515w4516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4523w4524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4531w4532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4539w4540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4547w4548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4555w4556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4411w4412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4563w4564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4571w4572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4579w4580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4587w4588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4595w4596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4603w4604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4611w4612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4619w4620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4627w4628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4635w4636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4419w4420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4643w4644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4651w4652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4427w4428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4435w4436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4443w4444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4451w4452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4459w4460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4467w4468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4475w4476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5178w5179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5259w5260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5267w5268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5275w5276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5283w5284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5291w5292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5299w5300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5307w5308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5315w5316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5323w5324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5331w5332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5187w5188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5339w5340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5347w5348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5355w5356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5363w5364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5371w5372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5379w5380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5387w5388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5395w5396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5403w5404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5411w5412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5195w5196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5419w5420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5427w5428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5203w5204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5211w5212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5219w5220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5227w5228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5235w5236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5243w5244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5251w5252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5949w5950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6030w6031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6038w6039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6046w6047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6054w6055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6062w6063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6070w6071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6078w6079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6086w6087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6094w6095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6102w6103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5958w5959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6110w6111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6118w6119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6126w6127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6134w6135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6142w6143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6150w6151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6158w6159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6166w6167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6174w6175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6182w6183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5966w5967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6190w6191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6198w6199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5974w5975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5982w5983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5990w5991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5998w5999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6006w6007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6014w6015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6022w6023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6715w6716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6796w6797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6804w6805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6812w6813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6820w6821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6828w6829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6836w6837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6844w6845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6852w6853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6860w6861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6868w6869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6724w6725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6876w6877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6884w6885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6892w6893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6900w6901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6908w6909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6916w6917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6924w6925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6932w6933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6940w6941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6948w6949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6732w6733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6956w6957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6964w6965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6740w6741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6748w6749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6756w6757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6764w6765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6772w6773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6780w6781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6788w6789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7476w7477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7557w7558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7565w7566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7573w7574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7581w7582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7589w7590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7597w7598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7605w7606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7613w7614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7621w7622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7629w7630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7485w7486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7637w7638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7645w7646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7653w7654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7661w7662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7669w7670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7677w7678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7685w7686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7693w7694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7701w7702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7709w7710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7493w7494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7717w7718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7725w7726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7501w7502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7509w7510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7517w7518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7525w7526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7533w7534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7541w7542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7549w7550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range9996w9997w9998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10033w10050w10051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10038w10055w10056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10043w10060w10061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10048w10065w10066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10053w10070w10071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10058w10075w10076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10063w10080w10081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10068w10085w10086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10073w10090w10091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10078w10095w10096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10003w10004w10005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10083w10100w10101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10088w10105w10106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10093w10110w10111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10098w10115w10116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10103w10120w10121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10108w10125w10126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10113w10130w10131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10118w10135w10136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10123w10140w10141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10128w10143w10144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10009w10010w10011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10133w10146w10147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10138w10149w10150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range9993w10015w10016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10001w10020w10021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10007w10025w10026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10013w10030w10031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10018w10035w10036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10023w10040w10041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10028w10045w10046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range335w338w339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range340w343w344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range345w348w349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range350w353w354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range355w358w359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range360w363w364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range365w368w369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range370w373w374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range375w378w379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range380w383w384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range385w388w389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range390w393w394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range395w398w399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range400w403w404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range405w408w409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range410w413w414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range415w418w419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range420w423w424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range425w428w429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range430w433w434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range435w438w439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range440w443w444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range300w303w304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range305w308w309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range310w313w314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range315w318w319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range320w323w324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range325w328w329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_radians_range330w333w334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7019w7212w7213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7078w7294w7295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7084w7302w7303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7090w7310w7311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7096w7318w7319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7102w7326w7327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7108w7334w7335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7114w7342w7343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7120w7350w7351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7126w7358w7359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7132w7366w7367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7024w7222w7223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7138w7374w7375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7144w7382w7383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7148w7390w7391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6970w7398w7399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6975w7406w7407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6977w7414w7415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6979w7422w7423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6981w7430w7431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6983w7438w7439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6985w7446w7447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7030w7230w7231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6987w7454w7455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6989w7462w7463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7036w7238w7239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7042w7246w7247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7048w7254w7255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7054w7262w7263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7060w7270w7271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7066w7278w7279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7072w7286w7287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7784w7968w7969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7843w8050w8051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7849w8058w8059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7855w8066w8067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7861w8074w8075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7867w8082w8083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7873w8090w8091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7879w8098w8099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7885w8106w8107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7891w8114w8115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7897w8122w8123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7789w7978w7979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7903w8130w8131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7907w8138w8139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7731w8146w8147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7736w8154w8155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7738w8162w8163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7740w8170w8171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7742w8178w8179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7744w8186w8187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7746w8194w8195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7748w8202w8203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7795w7986w7987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7750w8210w8211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7752w8218w8219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7801w7994w7995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7807w8002w8003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7813w8010w8011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7819w8018w8019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7825w8026w8027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7831w8034w8035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7837w8042w8043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8544w8719w8720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8603w8801w8802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8609w8809w8810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8615w8817w8818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8621w8825w8826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8627w8833w8834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8633w8841w8842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8639w8849w8850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8645w8857w8858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8651w8865w8866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8657w8873w8874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8549w8729w8730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8661w8881w8882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8487w8889w8890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8492w8897w8898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8494w8905w8906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8496w8913w8914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8498w8921w8922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8500w8929w8930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8502w8937w8938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8504w8945w8946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8506w8953w8954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8555w8737w8738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8508w8961w8962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8510w8969w8970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8561w8745w8746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8567w8753w8754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8573w8761w8762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8579w8769w8770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8585w8777w8778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8591w8785w8786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8597w8793w8794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9299w9465w9466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9358w9547w9548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9364w9555w9556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9370w9563w9564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9376w9571w9572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9382w9579w9580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9388w9587w9588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9394w9595w9596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9400w9603w9604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9406w9611w9612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9410w9619w9620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9304w9475w9476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9238w9627w9628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9243w9635w9636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9245w9643w9644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9247w9651w9652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9249w9659w9660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9251w9667w9668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9253w9675w9676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9255w9683w9684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9257w9691w9692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9259w9699w9700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9310w9483w9484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9261w9707w9708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9263w9715w9716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9316w9491w9492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9322w9499w9500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9328w9507w9508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9334w9515w9516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9340w9523w9524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9346w9531w9532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9352w9539w9540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range719w984w985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range778w1066w1067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range784w1074w1075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range790w1082w1083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range796w1090w1091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range802w1098w1099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range808w1106w1107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range814w1114w1115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range820w1122w1123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range826w1130w1131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range832w1138w1139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range724w994w995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range838w1146w1147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range844w1154w1155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range850w1162w1163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range856w1170w1171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range862w1178w1179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range868w1186w1187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range874w1194w1195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range880w1202w1203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range886w1210w1211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range892w1218w1219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range730w1002w1003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range896w1226w1227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range702w1234w1235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range736w1010w1011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range742w1018w1019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range748w1026w1027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range754w1034w1035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range760w1042w1043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range766w1050w1051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range772w1058w1059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1524w1780w1781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1583w1862w1863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1589w1870w1871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1595w1878w1879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1601w1886w1887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1607w1894w1895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1613w1902w1903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1619w1910w1911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1625w1918w1919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1631w1926w1927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1637w1934w1935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1529w1790w1791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1643w1942w1943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1649w1950w1951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1655w1958w1959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1661w1966w1967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1667w1974w1975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1673w1982w1983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1679w1990w1991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1685w1998w1999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1691w2006w2007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1695w2014w2015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1535w1798w1799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1503w2022w2023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1508w2030w2031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1541w1806w1807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1547w1814w1815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1553w1822w1823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1559w1830w1831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1565w1838w1839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1571w1846w1847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1577w1854w1855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2324w2571w2572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2383w2653w2654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2389w2661w2662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2395w2669w2670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2401w2677w2678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2407w2685w2686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2413w2693w2694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2419w2701w2702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2425w2709w2710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2431w2717w2718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2437w2725w2726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2329w2581w2582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2443w2733w2734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2449w2741w2742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2455w2749w2750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2461w2757w2758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2467w2765w2766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2473w2773w2774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2479w2781w2782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2485w2789w2790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2489w2797w2798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2299w2805w2806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2335w2589w2590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2304w2813w2814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2306w2821w2822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2341w2597w2598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2347w2605w2606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2353w2613w2614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2359w2621w2622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2365w2629w2630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2371w2637w2638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2377w2645w2646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3119w3357w3358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3178w3439w3440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3184w3447w3448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3190w3455w3456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3196w3463w3464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3202w3471w3472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3208w3479w3480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3214w3487w3488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3220w3495w3496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3226w3503w3504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3232w3511w3512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3124w3367w3368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3238w3519w3520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3244w3527w3528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3250w3535w3536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3256w3543w3544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3262w3551w3552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3268w3559w3560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3274w3567w3568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3278w3575w3576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3090w3583w3584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3095w3591w3592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3130w3375w3376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3097w3599w3600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3099w3607w3608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3136w3383w3384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3142w3391w3392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3148w3399w3400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3154w3407w3408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3160w3415w3416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3166w3423w3424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3172w3431w3432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3909w4138w4139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3968w4220w4221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3974w4228w4229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3980w4236w4237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3986w4244w4245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3992w4252w4253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3998w4260w4261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4004w4268w4269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4010w4276w4277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4016w4284w4285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4022w4292w4293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3914w4148w4149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4028w4300w4301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4034w4308w4309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4040w4316w4317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4046w4324w4325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4052w4332w4333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4058w4340w4341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4062w4348w4349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3876w4356w4357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3881w4364w4365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3883w4372w4373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3920w4156w4157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3885w4380w4381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3887w4388w4389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3926w4164w4165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3932w4172w4173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3938w4180w4181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3944w4188w4189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3950w4196w4197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3956w4204w4205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3962w4212w4213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4694w4914w4915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4753w4996w4997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4759w5004w5005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4765w5012w5013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4771w5020w5021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4777w5028w5029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4783w5036w5037w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4789w5044w5045w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4795w5052w5053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4801w5060w5061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4807w5068w5069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4699w4924w4925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4813w5076w5077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4819w5084w5085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4825w5092w5093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4831w5100w5101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4837w5108w5109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4841w5116w5117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4657w5124w5125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4662w5132w5133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4664w5140w5141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4666w5148w5149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4705w4932w4933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4668w5156w5157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4670w5164w5165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4711w4940w4941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4717w4948w4949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4723w4956w4957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4729w4964w4965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4735w4972w4973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4741w4980w4981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4747w4988w4989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5474w5685w5686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5533w5767w5768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5539w5775w5776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5545w5783w5784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5551w5791w5792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5557w5799w5800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5563w5807w5808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5569w5815w5816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5575w5823w5824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5581w5831w5832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5587w5839w5840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5479w5695w5696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5593w5847w5848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5599w5855w5856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5605w5863w5864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5611w5871w5872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5615w5879w5880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5433w5887w5888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5438w5895w5896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5440w5903w5904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5442w5911w5912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5444w5919w5920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5485w5703w5704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5446w5927w5928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5448w5935w5936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5491w5711w5712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5497w5719w5720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5503w5727w5728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5509w5735w5736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5515w5743w5744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5521w5751w5752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5527w5759w5760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6249w6451w6452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6308w6533w6534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6314w6541w6542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6320w6549w6550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6326w6557w6558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6332w6565w6566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6338w6573w6574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6344w6581w6582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6350w6589w6590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6356w6597w6598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6362w6605w6606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6254w6461w6462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6368w6613w6614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6374w6621w6622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6380w6629w6630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6384w6637w6638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6204w6645w6646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6209w6653w6654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6211w6661w6662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6213w6669w6670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6215w6677w6678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6217w6685w6686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6260w6469w6470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6219w6693w6694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6221w6701w6702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6266w6477w6478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6272w6485w6486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6278w6493w6494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6284w6501w6502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6290w6509w6510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6296w6517w6518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6302w6525w6526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7021w7217w7218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7080w7298w7299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7086w7306w7307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7092w7314w7315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7098w7322w7323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7104w7330w7331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7110w7338w7339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7116w7346w7347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7122w7354w7355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7128w7362w7363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7134w7370w7371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7026w7226w7227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7140w7378w7379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7146w7386w7387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7149w7394w7395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6973w7402w7403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6976w7410w7411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6978w7418w7419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6980w7426w7427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6982w7434w7435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6984w7442w7443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6986w7450w7451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7032w7234w7235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6988w7458w7459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6990w7466w7467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7038w7242w7243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7044w7250w7251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7050w7258w7259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7056w7266w7267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7062w7274w7275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7068w7282w7283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7074w7290w7291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7786w7973w7974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7845w8054w8055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7851w8062w8063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7857w8070w8071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7863w8078w8079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7869w8086w8087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7875w8094w8095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7881w8102w8103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7887w8110w8111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7893w8118w8119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7899w8126w8127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7791w7982w7983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7905w8134w8135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7908w8142w8143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7734w8150w8151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7737w8158w8159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7739w8166w8167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7741w8174w8175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7743w8182w8183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7745w8190w8191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7747w8198w8199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7749w8206w8207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7797w7990w7991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7751w8214w8215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7753w8222w8223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7803w7998w7999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7809w8006w8007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7815w8014w8015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7821w8022w8023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7827w8030w8031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7833w8038w8039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7839w8046w8047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8546w8724w8725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8605w8805w8806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8611w8813w8814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8617w8821w8822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8623w8829w8830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8629w8837w8838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8635w8845w8846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8641w8853w8854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8647w8861w8862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8653w8869w8870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8659w8877w8878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8551w8733w8734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8662w8885w8886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8490w8893w8894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8493w8901w8902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8495w8909w8910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8497w8917w8918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8499w8925w8926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8501w8933w8934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8503w8941w8942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8505w8949w8950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8507w8957w8958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8557w8741w8742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8509w8965w8966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8511w8973w8974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8563w8749w8750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8569w8757w8758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8575w8765w8766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8581w8773w8774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8587w8781w8782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8593w8789w8790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8599w8797w8798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9301w9470w9471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9360w9551w9552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9366w9559w9560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9372w9567w9568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9378w9575w9576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9384w9583w9584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9390w9591w9592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9396w9599w9600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9402w9607w9608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9408w9615w9616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9411w9623w9624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9306w9479w9480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9241w9631w9632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9244w9639w9640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9246w9647w9648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9248w9655w9656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9250w9663w9664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9252w9671w9672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9254w9679w9680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9256w9687w9688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9258w9695w9696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9260w9703w9704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9312w9487w9488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9262w9711w9712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9264w9719w9720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9318w9495w9496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9324w9503w9504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9330w9511w9512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9336w9519w9520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9342w9527w9528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9348w9535w9536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9354w9543w9544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range721w989w990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range780w1070w1071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range786w1078w1079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range792w1086w1087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range798w1094w1095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range804w1102w1103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range810w1110w1111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range816w1118w1119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range822w1126w1127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range828w1134w1135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range834w1142w1143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range726w998w999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range840w1150w1151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range846w1158w1159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range852w1166w1167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range858w1174w1175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range864w1182w1183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range870w1190w1191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range876w1198w1199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range882w1206w1207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range888w1214w1215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range894w1222w1223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range732w1006w1007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range897w1230w1231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range705w1238w1239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range738w1014w1015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range744w1022w1023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range750w1030w1031w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range756w1038w1039w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range762w1046w1047w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range768w1054w1055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range774w1062w1063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1526w1785w1786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1585w1866w1867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1591w1874w1875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1597w1882w1883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1603w1890w1891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1609w1898w1899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1615w1906w1907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1621w1914w1915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1627w1922w1923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1633w1930w1931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1639w1938w1939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1531w1794w1795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1645w1946w1947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1651w1954w1955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1657w1962w1963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1663w1970w1971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1669w1978w1979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1675w1986w1987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1681w1994w1995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1687w2002w2003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1693w2010w2011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1696w2018w2019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1537w1802w1803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1506w2026w2027w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1509w2034w2035w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1543w1810w1811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1549w1818w1819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1555w1826w1827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1561w1834w1835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1567w1842w1843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1573w1850w1851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1579w1858w1859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2326w2576w2577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2385w2657w2658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2391w2665w2666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2397w2673w2674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2403w2681w2682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2409w2689w2690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2415w2697w2698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2421w2705w2706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2427w2713w2714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2433w2721w2722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2439w2729w2730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2331w2585w2586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2445w2737w2738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2451w2745w2746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2457w2753w2754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2463w2761w2762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2469w2769w2770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2475w2777w2778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2481w2785w2786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2487w2793w2794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2490w2801w2802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2302w2809w2810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2337w2593w2594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2305w2817w2818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2307w2825w2826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2343w2601w2602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2349w2609w2610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2355w2617w2618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2361w2625w2626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2367w2633w2634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2373w2641w2642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2379w2649w2650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3121w3362w3363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3180w3443w3444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3186w3451w3452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3192w3459w3460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3198w3467w3468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3204w3475w3476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3210w3483w3484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3216w3491w3492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3222w3499w3500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3228w3507w3508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3234w3515w3516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3126w3371w3372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3240w3523w3524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3246w3531w3532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3252w3539w3540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3258w3547w3548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3264w3555w3556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3270w3563w3564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3276w3571w3572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3279w3579w3580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3093w3587w3588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3096w3595w3596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3132w3379w3380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3098w3603w3604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3100w3611w3612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3138w3387w3388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3144w3395w3396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3150w3403w3404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3156w3411w3412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3162w3419w3420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3168w3427w3428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3174w3435w3436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3911w4143w4144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3970w4224w4225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3976w4232w4233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3982w4240w4241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3988w4248w4249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3994w4256w4257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4000w4264w4265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4006w4272w4273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4012w4280w4281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4018w4288w4289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4024w4296w4297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3916w4152w4153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4030w4304w4305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4036w4312w4313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4042w4320w4321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4048w4328w4329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4054w4336w4337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4060w4344w4345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4063w4352w4353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3879w4360w4361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3882w4368w4369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3884w4376w4377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3922w4160w4161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3886w4384w4385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3888w4392w4393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3928w4168w4169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3934w4176w4177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3940w4184w4185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3946w4192w4193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3952w4200w4201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3958w4208w4209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3964w4216w4217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4696w4919w4920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4755w5000w5001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4761w5008w5009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4767w5016w5017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4773w5024w5025w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4779w5032w5033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4785w5040w5041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4791w5048w5049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4797w5056w5057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4803w5064w5065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4809w5072w5073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4701w4928w4929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4815w5080w5081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4821w5088w5089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4827w5096w5097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4833w5104w5105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4839w5112w5113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4842w5120w5121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4660w5128w5129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4663w5136w5137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4665w5144w5145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4667w5152w5153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4707w4936w4937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4669w5160w5161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4671w5168w5169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4713w4944w4945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4719w4952w4953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4725w4960w4961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4731w4968w4969w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4737w4976w4977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4743w4984w4985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4749w4992w4993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5476w5690w5691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5535w5771w5772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5541w5779w5780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5547w5787w5788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5553w5795w5796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5559w5803w5804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5565w5811w5812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5571w5819w5820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5577w5827w5828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5583w5835w5836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5589w5843w5844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5481w5699w5700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5595w5851w5852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5601w5859w5860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5607w5867w5868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5613w5875w5876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5616w5883w5884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5436w5891w5892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5439w5899w5900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5441w5907w5908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5443w5915w5916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5445w5923w5924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5487w5707w5708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5447w5931w5932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5449w5939w5940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5493w5715w5716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5499w5723w5724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5505w5731w5732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5511w5739w5740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5517w5747w5748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5523w5755w5756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5529w5763w5764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6251w6456w6457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6310w6537w6538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6316w6545w6546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6322w6553w6554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6328w6561w6562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6334w6569w6570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6340w6577w6578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6346w6585w6586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6352w6593w6594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6358w6601w6602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6364w6609w6610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6256w6465w6466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6370w6617w6618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6376w6625w6626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6382w6633w6634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6385w6641w6642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6207w6649w6650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6210w6657w6658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6212w6665w6666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6214w6673w6674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6216w6681w6682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6218w6689w6690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6262w6473w6474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6220w6697w6698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6222w6705w6706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6268w6481w6482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6274w6489w6490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6280w6497w6498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6286w6505w6506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6292w6513w6514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6298w6521w6522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6304w6529w6530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8232w8233w8234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8313w8314w8315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8321w8322w8323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8329w8330w8331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8337w8338w8339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8345w8346w8347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8353w8354w8355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8361w8362w8363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8369w8370w8371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8377w8378w8379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8385w8386w8387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8241w8242w8243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8393w8394w8395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8401w8402w8403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8409w8410w8411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8417w8418w8419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8425w8426w8427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8433w8434w8435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8441w8442w8443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8449w8450w8451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8457w8458w8459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8465w8466w8467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8249w8250w8251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8473w8474w8475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8481w8482w8483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8257w8258w8259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8265w8266w8267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8273w8274w8275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8281w8282w8283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8289w8290w8291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8297w8298w8299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8305w8306w8307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range8983w8984w8985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9064w9065w9066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9072w9073w9074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9080w9081w9082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9088w9089w9090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9096w9097w9098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9104w9105w9106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9112w9113w9114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9120w9121w9122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9128w9129w9130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9136w9137w9138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range8992w8993w8994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9144w9145w9146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9152w9153w9154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9160w9161w9162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9168w9169w9170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9176w9177w9178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9184w9185w9186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9192w9193w9194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9200w9201w9202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9208w9209w9210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9216w9217w9218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9000w9001w9002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9224w9225w9226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9232w9233w9234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9008w9009w9010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9016w9017w9018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9024w9025w9026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9032w9033w9034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9040w9041w9042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9048w9049w9050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9056w9057w9058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9729w9730w9731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9810w9811w9812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9818w9819w9820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9826w9827w9828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9834w9835w9836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9842w9843w9844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9850w9851w9852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9858w9859w9860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9866w9867w9868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9874w9875w9876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9882w9883w9884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9738w9739w9740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9890w9891w9892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9898w9899w9900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9906w9907w9908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9914w9915w9916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9922w9923w9924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9930w9931w9932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9938w9939w9940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9946w9947w9948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9954w9955w9956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9962w9963w9964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9746w9747w9748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9970w9971w9972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9978w9979w9980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9754w9755w9756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9762w9763w9764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9770w9771w9772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9778w9779w9780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9786w9787w9788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9794w9795w9796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9802w9803w9804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1248w1249w1250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1329w1330w1331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1337w1338w1339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1345w1346w1347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1353w1354w1355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1361w1362w1363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1369w1370w1371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1377w1378w1379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1385w1386w1387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1393w1394w1395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1401w1402w1403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1257w1258w1259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1409w1410w1411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1417w1418w1419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1425w1426w1427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1433w1434w1435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1441w1442w1443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1449w1450w1451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1457w1458w1459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1465w1466w1467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1473w1474w1475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1481w1482w1483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1265w1266w1267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1489w1490w1491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1497w1498w1499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1273w1274w1275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1281w1282w1283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1289w1290w1291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1297w1298w1299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1305w1306w1307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1313w1314w1315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1321w1322w1323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2044w2045w2046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2125w2126w2127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2133w2134w2135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2141w2142w2143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2149w2150w2151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2157w2158w2159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2165w2166w2167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2173w2174w2175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2181w2182w2183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2189w2190w2191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2197w2198w2199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2053w2054w2055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2205w2206w2207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2213w2214w2215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2221w2222w2223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2229w2230w2231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2237w2238w2239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2245w2246w2247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2253w2254w2255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2261w2262w2263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2269w2270w2271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2277w2278w2279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2061w2062w2063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2285w2286w2287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2293w2294w2295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2069w2070w2071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2077w2078w2079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2085w2086w2087w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2093w2094w2095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2101w2102w2103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2109w2110w2111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2117w2118w2119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2835w2836w2837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2916w2917w2918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2924w2925w2926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2932w2933w2934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2940w2941w2942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2948w2949w2950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2956w2957w2958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2964w2965w2966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2972w2973w2974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2980w2981w2982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2988w2989w2990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2844w2845w2846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2996w2997w2998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3004w3005w3006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3012w3013w3014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3020w3021w3022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3028w3029w3030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3036w3037w3038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3044w3045w3046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3052w3053w3054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3060w3061w3062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3068w3069w3070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2852w2853w2854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3076w3077w3078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3084w3085w3086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2860w2861w2862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2868w2869w2870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2876w2877w2878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2884w2885w2886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2892w2893w2894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2900w2901w2902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2908w2909w2910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3621w3622w3623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3702w3703w3704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3710w3711w3712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3718w3719w3720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3726w3727w3728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3734w3735w3736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3742w3743w3744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3750w3751w3752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3758w3759w3760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3766w3767w3768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3774w3775w3776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3630w3631w3632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3782w3783w3784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3790w3791w3792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3798w3799w3800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3806w3807w3808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3814w3815w3816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3822w3823w3824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3830w3831w3832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3838w3839w3840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3846w3847w3848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3854w3855w3856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3638w3639w3640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3862w3863w3864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3870w3871w3872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3646w3647w3648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3654w3655w3656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3662w3663w3664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3670w3671w3672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3678w3679w3680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3686w3687w3688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3694w3695w3696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4402w4403w4404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4483w4484w4485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4491w4492w4493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4499w4500w4501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4507w4508w4509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4515w4516w4517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4523w4524w4525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4531w4532w4533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4539w4540w4541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4547w4548w4549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4555w4556w4557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4411w4412w4413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4563w4564w4565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4571w4572w4573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4579w4580w4581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4587w4588w4589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4595w4596w4597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4603w4604w4605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4611w4612w4613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4619w4620w4621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4627w4628w4629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4635w4636w4637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4419w4420w4421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4643w4644w4645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4651w4652w4653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4427w4428w4429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4435w4436w4437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4443w4444w4445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4451w4452w4453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4459w4460w4461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4467w4468w4469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4475w4476w4477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5178w5179w5180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5259w5260w5261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5267w5268w5269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5275w5276w5277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5283w5284w5285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5291w5292w5293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5299w5300w5301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5307w5308w5309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5315w5316w5317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5323w5324w5325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5331w5332w5333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5187w5188w5189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5339w5340w5341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5347w5348w5349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5355w5356w5357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5363w5364w5365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5371w5372w5373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5379w5380w5381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5387w5388w5389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5395w5396w5397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5403w5404w5405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5411w5412w5413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5195w5196w5197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5419w5420w5421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5427w5428w5429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5203w5204w5205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5211w5212w5213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5219w5220w5221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5227w5228w5229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5235w5236w5237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5243w5244w5245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5251w5252w5253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5949w5950w5951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6030w6031w6032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6038w6039w6040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6046w6047w6048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6054w6055w6056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6062w6063w6064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6070w6071w6072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6078w6079w6080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6086w6087w6088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6094w6095w6096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6102w6103w6104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5958w5959w5960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6110w6111w6112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6118w6119w6120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6126w6127w6128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6134w6135w6136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6142w6143w6144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6150w6151w6152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6158w6159w6160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6166w6167w6168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6174w6175w6176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6182w6183w6184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5966w5967w5968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6190w6191w6192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6198w6199w6200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5974w5975w5976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5982w5983w5984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5990w5991w5992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5998w5999w6000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6006w6007w6008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6014w6015w6016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6022w6023w6024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6715w6716w6717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6796w6797w6798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6804w6805w6806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6812w6813w6814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6820w6821w6822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6828w6829w6830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6836w6837w6838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6844w6845w6846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6852w6853w6854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6860w6861w6862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6868w6869w6870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6724w6725w6726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6876w6877w6878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6884w6885w6886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6892w6893w6894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6900w6901w6902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6908w6909w6910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6916w6917w6918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6924w6925w6926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6932w6933w6934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6940w6941w6942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6948w6949w6950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6732w6733w6734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6956w6957w6958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6964w6965w6966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6740w6741w6742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6748w6749w6750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6756w6757w6758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6764w6765w6766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6772w6773w6774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6780w6781w6782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6788w6789w6790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7476w7477w7478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7557w7558w7559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7565w7566w7567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7573w7574w7575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7581w7582w7583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7589w7590w7591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7597w7598w7599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7605w7606w7607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7613w7614w7615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7621w7622w7623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7629w7630w7631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7485w7486w7487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7637w7638w7639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7645w7646w7647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7653w7654w7655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7661w7662w7663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7669w7670w7671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7677w7678w7679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7685w7686w7687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7693w7694w7695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7701w7702w7703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7709w7710w7711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7493w7494w7495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7717w7718w7719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7725w7726w7727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7501w7502w7503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7509w7510w7511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7517w7518w7519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7525w7526w7527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7533w7534w7535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7541w7542w7543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7549w7550w7551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_estimate_w10152w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7214w7470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7296w7553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7304w7561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7312w7569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7320w7577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7328w7585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7336w7593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7344w7601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7352w7609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7360w7617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7368w7625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7224w7481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7376w7633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7384w7641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7392w7649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7400w7657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7408w7665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7416w7673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7424w7681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7432w7689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7440w7697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7448w7705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7232w7489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7456w7713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7464w7721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7240w7497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7248w7505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7256w7513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7264w7521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7272w7529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7280w7537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7288w7545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range7970w8226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8052w8309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8060w8317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8068w8325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8076w8333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8084w8341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8092w8349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8100w8357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8108w8365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8116w8373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8124w8381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range7980w8237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8132w8389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8140w8397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8148w8405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8156w8413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8164w8421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8172w8429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8180w8437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8188w8445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8196w8453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8204w8461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range7988w8245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8212w8469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8220w8477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range7996w8253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8004w8261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8012w8269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8020w8277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8028w8285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8036w8293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8044w8301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8721w8977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8803w9060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8811w9068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8819w9076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8827w9084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8835w9092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8843w9100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8851w9108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8859w9116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8867w9124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8875w9132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8731w8988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8883w9140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8891w9148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8899w9156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8907w9164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8915w9172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8923w9180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8931w9188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8939w9196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8947w9204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8955w9212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8739w8996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8963w9220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8971w9228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8747w9004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8755w9012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8763w9020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8771w9028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8779w9036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8787w9044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8795w9052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9467w9723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9549w9806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9557w9814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9565w9822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9573w9830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9581w9838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9589w9846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9597w9854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9605w9862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9613w9870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9621w9878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9477w9734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9629w9886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9637w9894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9645w9902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9653w9910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9661w9918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9669w9926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9677w9934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9685w9942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9693w9950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9701w9958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9485w9742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9709w9966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9717w9974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9493w9750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9501w9758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9509w9766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9517w9774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9525w9782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9533w9790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9541w9798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range986w1242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1068w1325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1076w1333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1084w1341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1092w1349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1100w1357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1108w1365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1116w1373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1124w1381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1132w1389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1140w1397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range996w1253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1148w1405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1156w1413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1164w1421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1172w1429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1180w1437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1188w1445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1196w1453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1204w1461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1212w1469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1220w1477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1004w1261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1228w1485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1236w1493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1012w1269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1020w1277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1028w1285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1036w1293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1044w1301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1052w1309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1060w1317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1782w2038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1864w2121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1872w2129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1880w2137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1888w2145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1896w2153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1904w2161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1912w2169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1920w2177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1928w2185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1936w2193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1792w2049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1944w2201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1952w2209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1960w2217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1968w2225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1976w2233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1984w2241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1992w2249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2000w2257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2008w2265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2016w2273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1800w2057w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2024w2281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2032w2289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1808w2065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1816w2073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1824w2081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1832w2089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1840w2097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1848w2105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1856w2113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2573w2829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2655w2912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2663w2920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2671w2928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2679w2936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2687w2944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2695w2952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2703w2960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2711w2968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2719w2976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2727w2984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2583w2840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2735w2992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2743w3000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2751w3008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2759w3016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2767w3024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2775w3032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2783w3040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2791w3048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2799w3056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2807w3064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2591w2848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2815w3072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2823w3080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2599w2856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2607w2864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2615w2872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2623w2880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2631w2888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2639w2896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2647w2904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3359w3615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3441w3698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3449w3706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3457w3714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3465w3722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3473w3730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3481w3738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3489w3746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3497w3754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3505w3762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3513w3770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3369w3626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3521w3778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3529w3786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3537w3794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3545w3802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3553w3810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3561w3818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3569w3826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3577w3834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3585w3842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3593w3850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3377w3634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3601w3858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3609w3866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3385w3642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3393w3650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3401w3658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3409w3666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3417w3674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3425w3682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3433w3690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4140w4396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4222w4479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4230w4487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4238w4495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4246w4503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4254w4511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4262w4519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4270w4527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4278w4535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4286w4543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4294w4551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4150w4407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4302w4559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4310w4567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4318w4575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4326w4583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4334w4591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4342w4599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4350w4607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4358w4615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4366w4623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4374w4631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4158w4415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4382w4639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4390w4647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4166w4423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4174w4431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4182w4439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4190w4447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4198w4455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4206w4463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4214w4471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4916w5172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4998w5255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5006w5263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5014w5271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5022w5279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5030w5287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5038w5295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5046w5303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5054w5311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5062w5319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5070w5327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4926w5183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5078w5335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5086w5343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5094w5351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5102w5359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5110w5367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5118w5375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5126w5383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5134w5391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5142w5399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5150w5407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4934w5191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5158w5415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5166w5423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4942w5199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4950w5207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4958w5215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4966w5223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4974w5231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4982w5239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4990w5247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5687w5943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5769w6026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5777w6034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5785w6042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5793w6050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5801w6058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5809w6066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5817w6074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5825w6082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5833w6090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5841w6098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5697w5954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5849w6106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5857w6114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5865w6122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5873w6130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5881w6138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5889w6146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5897w6154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5905w6162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5913w6170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5921w6178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5705w5962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5929w6186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5937w6194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5713w5970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5721w5978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5729w5986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5737w5994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5745w6002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5753w6010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5761w6018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6453w6709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6535w6792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6543w6800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6551w6808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6559w6816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6567w6824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6575w6832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6583w6840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6591w6848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6599w6856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6607w6864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6463w6720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6615w6872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6623w6880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6631w6888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6639w6896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6647w6904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6655w6912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6663w6920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6671w6928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6679w6936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6687w6944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6471w6728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6695w6952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6703w6960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6479w6736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6487w6744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6495w6752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6503w6760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6511w6768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6519w6776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6527w6784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7219w7473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7300w7555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7308w7563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7316w7571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7324w7579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7332w7587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7340w7595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7348w7603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7356w7611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7364w7619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7372w7627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7228w7483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7380w7635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7388w7643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7396w7651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7404w7659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7412w7667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7420w7675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7428w7683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7436w7691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7444w7699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7452w7707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7236w7491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7460w7715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7468w7723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7244w7499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7252w7507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7260w7515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7268w7523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7276w7531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7284w7539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7292w7547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range7975w8229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8056w8311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8064w8319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8072w8327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8080w8335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8088w8343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8096w8351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8104w8359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8112w8367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8120w8375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8128w8383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range7984w8239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8136w8391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8144w8399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8152w8407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8160w8415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8168w8423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8176w8431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8184w8439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8192w8447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8200w8455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8208w8463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range7992w8247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8216w8471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8224w8479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8000w8255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8008w8263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8016w8271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8024w8279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8032w8287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8040w8295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8048w8303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8726w8980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8807w9062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8815w9070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8823w9078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8831w9086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8839w9094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8847w9102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8855w9110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8863w9118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8871w9126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8879w9134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8735w8990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8887w9142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8895w9150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8903w9158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8911w9166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8919w9174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8927w9182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8935w9190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8943w9198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8951w9206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8959w9214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8743w8998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8967w9222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8975w9230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8751w9006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8759w9014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8767w9022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8775w9030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8783w9038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8791w9046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8799w9054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9472w9726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9553w9808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9561w9816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9569w9824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9577w9832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9585w9840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9593w9848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9601w9856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9609w9864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9617w9872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9625w9880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9481w9736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9633w9888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9641w9896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9649w9904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9657w9912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9665w9920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9673w9928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9681w9936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9689w9944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9697w9952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9705w9960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9489w9744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9713w9968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9721w9976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9497w9752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9505w9760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9513w9768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9521w9776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9529w9784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9537w9792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9545w9800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range991w1245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1072w1327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1080w1335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1088w1343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1096w1351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1104w1359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1112w1367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1120w1375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1128w1383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1136w1391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1144w1399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1000w1255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1152w1407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1160w1415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1168w1423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1176w1431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1184w1439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1192w1447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1200w1455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1208w1463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1216w1471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1224w1479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1008w1263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1232w1487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1240w1495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1016w1271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1024w1279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1032w1287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1040w1295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1048w1303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1056w1311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1064w1319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1787w2041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1868w2123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1876w2131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1884w2139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1892w2147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1900w2155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1908w2163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1916w2171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1924w2179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1932w2187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1940w2195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1796w2051w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1948w2203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1956w2211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1964w2219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1972w2227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1980w2235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1988w2243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1996w2251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2004w2259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2012w2267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2020w2275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1804w2059w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2028w2283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2036w2291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1812w2067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1820w2075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1828w2083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1836w2091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1844w2099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1852w2107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1860w2115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2578w2832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2659w2914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2667w2922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2675w2930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2683w2938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2691w2946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2699w2954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2707w2962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2715w2970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2723w2978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2731w2986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2587w2842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2739w2994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2747w3002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2755w3010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2763w3018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2771w3026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2779w3034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2787w3042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2795w3050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2803w3058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2811w3066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2595w2850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2819w3074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2827w3082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2603w2858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2611w2866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2619w2874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2627w2882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2635w2890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2643w2898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2651w2906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3364w3618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3445w3700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3453w3708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3461w3716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3469w3724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3477w3732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3485w3740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3493w3748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3501w3756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3509w3764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3517w3772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3373w3628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3525w3780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3533w3788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3541w3796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3549w3804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3557w3812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3565w3820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3573w3828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3581w3836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3589w3844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3597w3852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3381w3636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3605w3860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3613w3868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3389w3644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3397w3652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3405w3660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3413w3668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3421w3676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3429w3684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3437w3692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4145w4399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4226w4481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4234w4489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4242w4497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4250w4505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4258w4513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4266w4521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4274w4529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4282w4537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4290w4545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4298w4553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4154w4409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4306w4561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4314w4569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4322w4577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4330w4585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4338w4593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4346w4601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4354w4609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4362w4617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4370w4625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4378w4633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4162w4417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4386w4641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4394w4649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4170w4425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4178w4433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4186w4441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4194w4449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4202w4457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4210w4465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4218w4473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4921w5175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5002w5257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5010w5265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5018w5273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5026w5281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5034w5289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5042w5297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5050w5305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5058w5313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5066w5321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5074w5329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4930w5185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5082w5337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5090w5345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5098w5353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5106w5361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5114w5369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5122w5377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5130w5385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5138w5393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5146w5401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5154w5409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4938w5193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5162w5417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5170w5425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4946w5201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4954w5209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4962w5217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4970w5225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4978w5233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4986w5241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4994w5249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5692w5946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5773w6028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5781w6036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5789w6044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5797w6052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5805w6060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5813w6068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5821w6076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5829w6084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5837w6092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5845w6100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5701w5956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5853w6108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5861w6116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5869w6124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5877w6132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5885w6140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5893w6148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5901w6156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5909w6164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5917w6172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5925w6180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5709w5964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5933w6188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5941w6196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5717w5972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5725w5980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5733w5988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5741w5996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5749w6004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5757w6012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5765w6020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6458w6712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6539w6794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6547w6802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6555w6810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6563w6818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6571w6826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6579w6834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6587w6842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6595w6850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6603w6858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6611w6866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6467w6722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6619w6874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6627w6882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6635w6890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6643w6898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6651w6906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6659w6914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6667w6922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6675w6930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6683w6938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6691w6946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6475w6730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6699w6954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6707w6962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6483w6738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6491w6746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6499w6754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6507w6762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6515w6770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6523w6778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6531w6786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  atannode_0_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  atannode_10_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  atannode_11_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  atannode_12_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  atannode_1_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  atannode_2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  atannode_3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  atannode_4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  atannode_5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  atannode_6_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  atannode_7_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  atannode_8_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  atannode_9_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  delay_input_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  delay_pipe_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  estimate_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  indexpointnum_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  multiplier_input_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  multipliernode_w :	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  post_estimate_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  pre_estimate_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  radians_load_node_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  startindex_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  x_pipenode_10_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_pipenode_11_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_pipenode_12_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_pipenode_13_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_pipenode_2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_pipenode_3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_pipenode_4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_pipenode_5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_pipenode_6_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_pipenode_7_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_pipenode_8_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_pipenode_9_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenode_10_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenode_11_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenode_12_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenode_13_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenode_2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenode_3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenode_4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenode_5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenode_6_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenode_7_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenode_8_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenode_9_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodeone_10_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodeone_11_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodeone_12_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodeone_13_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodeone_2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodeone_3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodeone_4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodeone_5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodeone_6_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodeone_7_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodeone_8_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodeone_9_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodetwo_10_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodetwo_11_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodetwo_12_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodetwo_13_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodetwo_2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodetwo_3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodetwo_4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodetwo_5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodetwo_6_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodetwo_7_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodetwo_8_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_prenodetwo_9_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_start_node_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_subnode_10_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_subnode_11_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_subnode_12_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_subnode_13_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_subnode_2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_subnode_3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_subnode_4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_subnode_5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_subnode_6_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_subnode_7_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_subnode_8_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  x_subnode_9_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_pipenode_10_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_pipenode_11_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_pipenode_12_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_pipenode_13_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_pipenode_2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_pipenode_3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_pipenode_4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_pipenode_5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_pipenode_6_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_pipenode_7_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_pipenode_8_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_pipenode_9_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenode_10_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenode_11_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenode_12_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenode_13_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenode_2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenode_3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenode_4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenode_5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenode_6_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenode_7_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenode_8_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenode_9_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodeone_10_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodeone_11_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodeone_12_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodeone_13_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodeone_2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodeone_3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodeone_4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodeone_5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodeone_6_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodeone_7_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodeone_8_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodeone_9_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodetwo_10_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodetwo_11_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodetwo_12_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodetwo_13_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodetwo_2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodetwo_3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodetwo_4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodetwo_5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodetwo_6_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodetwo_7_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodetwo_8_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_prenodetwo_9_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_subnode_10_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_subnode_11_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_subnode_12_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_subnode_13_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_subnode_1_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_subnode_2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_subnode_3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_subnode_4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_subnode_5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_subnode_6_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_subnode_7_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_subnode_8_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  y_subnode_9_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_pipenode_10_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_pipenode_11_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_pipenode_12_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_pipenode_13_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_pipenode_2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_pipenode_3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_pipenode_4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_pipenode_5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_pipenode_6_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_pipenode_7_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_pipenode_8_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_pipenode_9_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_subnode_10_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_subnode_11_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_subnode_12_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_subnode_13_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_subnode_2_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_subnode_3_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_subnode_4_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_subnode_5_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_subnode_6_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_subnode_7_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_subnode_8_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  z_subnode_9_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_10_w_range8305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range8983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range8992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_11_w_range9056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9818w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9890w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_12_w_range9802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_1_w_range1321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2061w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2069w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_2_w_range2117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range3084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_3_w_range2908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3830w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_4_w_range3694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_5_w_range4475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_6_w_range5251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range5949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range5958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range5966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range5974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range5982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range5990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range5998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_7_w_range6022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_8_w_range6788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_atannode_9_w_range7549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range9996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10053w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range9993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_pre_estimate_w_range10028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_radians_range330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_10_w_range7288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range7970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range7980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range7988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range7996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_11_w_range8044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_12_w_range8795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_13_w_range9541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_2_w_range1060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range2032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_3_w_range1856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_4_w_range2647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_5_w_range3433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_6_w_range4214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range4916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range4998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range4926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range4934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range5166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range4942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range4950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range4958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range4966w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range4974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range4982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_7_w_range4990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5793w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5817w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_8_w_range5761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenode_9_w_range6527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range6970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range6975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range6977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range6979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range6981w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range6983w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range6985w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range6987w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range6989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_10_w_range7072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_11_w_range7837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_12_w_range8597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_13_w_range9352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range790w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range802w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range808w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range814w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range832w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_2_w_range772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1637w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_3_w_range1577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_4_w_range2377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_5_w_range3172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4046w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range4062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_6_w_range3962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4825w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_7_w_range4747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_8_w_range5527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodeone_9_w_range6302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range6991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range6995w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range6997w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range6999w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7005w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7009w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7939w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7942w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7945w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7957w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7960w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7963w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7912w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7915w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7778w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7918w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7936w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range979w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_2_w_range925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4097w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4067w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4070w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4073w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_10_w_range7292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range7975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range7984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range7992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_11_w_range8048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8823w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8831w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8903w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8927w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8967w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8975w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_12_w_range8799w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_13_w_range9545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1072w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1088w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1040w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_2_w_range1064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1796w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1972w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2028w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range2036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1836w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_3_w_range1860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2811w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_4_w_range2651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_5_w_range3437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_6_w_range4218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range4921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range4930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5090w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range4938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range5170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range4946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range4954w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range4962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range4970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range4978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range4986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_7_w_range4994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5805w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5829w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5837w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5885w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5909w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_8_w_range5765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenode_9_w_range6531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7026w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range6973w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range6976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range6978w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range6980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range6982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range6984w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range6986w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7032w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range6988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range6990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7038w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7044w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7062w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_10_w_range7074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7881w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7887w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7893w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7899w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_11_w_range7839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8647w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8662w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_12_w_range8599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_13_w_range9354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range828w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range834w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_2_w_range774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1597w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_3_w_range1579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2427w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_4_w_range2379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_5_w_range3174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3970w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3976w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3982w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3988w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3994w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4036w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4048w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4060w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range4063w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3882w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3888w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_6_w_range3964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4827w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4833w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_7_w_range4749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_8_w_range5529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6322w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodeone_9_w_range6304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range6993w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range6996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range6998w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7002w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7006w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7008w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7016w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7940w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7946w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7949w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7955w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7958w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7961w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7964w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7913w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7916w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7922w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7925w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7937w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8667w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8527w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9422w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range929w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range932w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range941w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range944w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range950w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range953w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range956w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range965w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range968w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range971w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range974w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range977w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range980w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range905w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range908w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range914w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range917w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_2_w_range926w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1704w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3332w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4098w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3891w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3894w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3902w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4077w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4089w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4883w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4886w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4889w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4892w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4895w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4898w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4901w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4904w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4910w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4677w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4859w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5657w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5672w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5627w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6432w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  coshw_altfp_sincos_cordic_atan_35b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_atan_k6b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_atan_l6b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_atan_m6b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_atan_n6b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_atan_45b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_atan_55b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_atan_65b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_atan_75b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_atan_85b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_atan_95b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_atan_a5b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_atan_b5b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_atan_c5b
	 PORT
	 ( 
		arctan	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		indexbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_cordic_start_509
	 PORT
	 ( 
		index	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
		value	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop30 : FOR i IN 0 TO 3 GENERATE 
		wire_ccc_cordic_m_w_lg_indexpointnum_w288w(i) <= indexpointnum_w(i) AND indexbit;
	END GENERATE loop30;
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range9996w9997w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range9996w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10033w10050w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10033w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10033w10034w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10033w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10038w10055w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10038w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10038w10039w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10038w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10043w10060w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10043w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10043w10044w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10043w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10048w10065w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10048w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10048w10049w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10048w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10053w10070w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10053w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10053w10054w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10053w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10058w10075w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10058w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10058w10059w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10058w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10063w10080w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10063w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10063w10064w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10063w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10068w10085w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10068w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10068w10069w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10068w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10073w10090w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10073w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10073w10074w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10073w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10078w10095w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10078w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10078w10079w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10078w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10003w10004w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10003w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10083w10100w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10083w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10083w10084w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10083w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10088w10105w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10088w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10088w10089w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10088w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10093w10110w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10093w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10093w10094w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10093w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10098w10115w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10098w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10098w10099w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10098w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10103w10120w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10103w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10103w10104w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10103w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10108w10125w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10108w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10108w10109w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10108w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10113w10130w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10113w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10113w10114w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10113w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10118w10135w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10118w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10118w10119w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10118w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10123w10140w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10123w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10123w10124w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10123w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10128w10143w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10128w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10128w10129w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10128w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10009w10010w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10009w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10133w10146w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10133w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10133w10134w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10133w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10138w10149w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10138w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10138w10139w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10138w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range9993w10015w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range9993w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range9993w9994w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range9993w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10001w10020w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10001w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10001w10002w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10001w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10007w10025w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10007w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10007w10008w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10007w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10013w10030w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10013w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10013w10014w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10013w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10018w10035w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10018w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10018w10019w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10018w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10023w10040w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10023w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10023w10024w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10023w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10028w10045w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10028w(0) AND wire_indexbitff_w_lg_w_q_range9992w9995w(0);
	wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10028w10029w(0) <= wire_ccc_cordic_m_w_pre_estimate_w_range10028w(0) AND wire_indexbitff_w_q_range9992w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range289w292w(0) <= wire_ccc_cordic_m_w_radians_range289w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range289w302w(0) <= wire_ccc_cordic_m_w_radians_range289w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range335w338w(0) <= wire_ccc_cordic_m_w_radians_range335w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range335w352w(0) <= wire_ccc_cordic_m_w_radians_range335w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range340w343w(0) <= wire_ccc_cordic_m_w_radians_range340w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range340w357w(0) <= wire_ccc_cordic_m_w_radians_range340w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range345w348w(0) <= wire_ccc_cordic_m_w_radians_range345w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range345w362w(0) <= wire_ccc_cordic_m_w_radians_range345w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range350w353w(0) <= wire_ccc_cordic_m_w_radians_range350w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range350w367w(0) <= wire_ccc_cordic_m_w_radians_range350w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range355w358w(0) <= wire_ccc_cordic_m_w_radians_range355w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range355w372w(0) <= wire_ccc_cordic_m_w_radians_range355w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range360w363w(0) <= wire_ccc_cordic_m_w_radians_range360w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range360w377w(0) <= wire_ccc_cordic_m_w_radians_range360w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range365w368w(0) <= wire_ccc_cordic_m_w_radians_range365w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range365w382w(0) <= wire_ccc_cordic_m_w_radians_range365w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range370w373w(0) <= wire_ccc_cordic_m_w_radians_range370w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range370w387w(0) <= wire_ccc_cordic_m_w_radians_range370w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range375w378w(0) <= wire_ccc_cordic_m_w_radians_range375w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range375w392w(0) <= wire_ccc_cordic_m_w_radians_range375w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range380w383w(0) <= wire_ccc_cordic_m_w_radians_range380w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range380w397w(0) <= wire_ccc_cordic_m_w_radians_range380w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range294w296w(0) <= wire_ccc_cordic_m_w_radians_range294w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range294w307w(0) <= wire_ccc_cordic_m_w_radians_range294w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range385w388w(0) <= wire_ccc_cordic_m_w_radians_range385w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range385w402w(0) <= wire_ccc_cordic_m_w_radians_range385w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range390w393w(0) <= wire_ccc_cordic_m_w_radians_range390w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range390w407w(0) <= wire_ccc_cordic_m_w_radians_range390w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range395w398w(0) <= wire_ccc_cordic_m_w_radians_range395w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range395w412w(0) <= wire_ccc_cordic_m_w_radians_range395w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range400w403w(0) <= wire_ccc_cordic_m_w_radians_range400w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range400w417w(0) <= wire_ccc_cordic_m_w_radians_range400w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range405w408w(0) <= wire_ccc_cordic_m_w_radians_range405w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range405w422w(0) <= wire_ccc_cordic_m_w_radians_range405w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range410w413w(0) <= wire_ccc_cordic_m_w_radians_range410w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range410w427w(0) <= wire_ccc_cordic_m_w_radians_range410w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range415w418w(0) <= wire_ccc_cordic_m_w_radians_range415w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range415w432w(0) <= wire_ccc_cordic_m_w_radians_range415w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range420w423w(0) <= wire_ccc_cordic_m_w_radians_range420w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range420w437w(0) <= wire_ccc_cordic_m_w_radians_range420w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range425w428w(0) <= wire_ccc_cordic_m_w_radians_range425w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range425w442w(0) <= wire_ccc_cordic_m_w_radians_range425w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range430w433w(0) <= wire_ccc_cordic_m_w_radians_range430w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range297w299w(0) <= wire_ccc_cordic_m_w_radians_range297w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range297w312w(0) <= wire_ccc_cordic_m_w_radians_range297w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range435w438w(0) <= wire_ccc_cordic_m_w_radians_range435w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range440w443w(0) <= wire_ccc_cordic_m_w_radians_range440w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range300w303w(0) <= wire_ccc_cordic_m_w_radians_range300w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range300w317w(0) <= wire_ccc_cordic_m_w_radians_range300w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range305w308w(0) <= wire_ccc_cordic_m_w_radians_range305w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range305w322w(0) <= wire_ccc_cordic_m_w_radians_range305w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range310w313w(0) <= wire_ccc_cordic_m_w_radians_range310w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range310w327w(0) <= wire_ccc_cordic_m_w_radians_range310w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range315w318w(0) <= wire_ccc_cordic_m_w_radians_range315w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range315w332w(0) <= wire_ccc_cordic_m_w_radians_range315w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range320w323w(0) <= wire_ccc_cordic_m_w_radians_range320w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range320w337w(0) <= wire_ccc_cordic_m_w_radians_range320w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range325w328w(0) <= wire_ccc_cordic_m_w_radians_range325w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range325w342w(0) <= wire_ccc_cordic_m_w_radians_range325w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_radians_range330w333w(0) <= wire_ccc_cordic_m_w_radians_range330w(0) AND wire_ccc_cordic_m_w_lg_indexbit291w(0);
	wire_ccc_cordic_m_w_lg_w_radians_range330w347w(0) <= wire_ccc_cordic_m_w_radians_range330w(0) AND indexbit;
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7019w7212w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7019w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7078w7294w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7078w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7084w7302w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7084w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7090w7310w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7090w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7096w7318w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7096w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7102w7326w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7102w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7108w7334w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7108w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7114w7342w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7114w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7120w7350w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7120w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7126w7358w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7126w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7132w7366w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7132w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7024w7222w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7024w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7138w7374w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7138w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7144w7382w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7144w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7148w7390w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7148w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6970w7398w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range6970w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6975w7406w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range6975w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6977w7414w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range6977w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6979w7422w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range6979w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6981w7430w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range6981w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6983w7438w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range6983w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6985w7446w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range6985w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7030w7230w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7030w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6987w7454w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range6987w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6989w7462w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range6989w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7036w7238w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7036w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7042w7246w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7042w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7048w7254w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7048w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7054w7262w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7054w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7060w7270w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7060w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7066w7278w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7066w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7072w7286w(0) <= wire_ccc_cordic_m_w_x_prenodeone_10_w_range7072w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7784w7968w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7784w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7843w8050w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7843w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7849w8058w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7849w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7855w8066w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7855w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7861w8074w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7861w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7867w8082w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7867w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7873w8090w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7873w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7879w8098w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7879w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7885w8106w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7885w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7891w8114w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7891w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7897w8122w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7897w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7789w7978w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7789w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7903w8130w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7903w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7907w8138w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7907w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7731w8146w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7731w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7736w8154w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7736w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7738w8162w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7738w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7740w8170w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7740w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7742w8178w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7742w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7744w8186w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7744w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7746w8194w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7746w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7748w8202w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7748w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7795w7986w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7795w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7750w8210w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7750w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7752w8218w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7752w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7801w7994w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7801w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7807w8002w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7807w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7813w8010w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7813w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7819w8018w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7819w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7825w8026w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7825w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7831w8034w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7831w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7837w8042w(0) <= wire_ccc_cordic_m_w_x_prenodeone_11_w_range7837w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8544w8719w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8544w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8603w8801w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8603w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8609w8809w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8609w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8615w8817w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8615w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8621w8825w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8621w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8627w8833w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8627w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8633w8841w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8633w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8639w8849w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8639w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8645w8857w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8645w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8651w8865w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8651w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8657w8873w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8657w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8549w8729w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8549w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8661w8881w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8661w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8487w8889w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8487w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8492w8897w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8492w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8494w8905w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8494w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8496w8913w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8496w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8498w8921w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8498w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8500w8929w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8500w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8502w8937w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8502w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8504w8945w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8504w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8506w8953w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8506w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8555w8737w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8555w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8508w8961w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8508w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8510w8969w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8510w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8561w8745w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8561w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8567w8753w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8567w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8573w8761w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8573w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8579w8769w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8579w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8585w8777w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8585w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8591w8785w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8591w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8597w8793w(0) <= wire_ccc_cordic_m_w_x_prenodeone_12_w_range8597w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9299w9465w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9299w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9358w9547w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9358w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9364w9555w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9364w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9370w9563w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9370w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9376w9571w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9376w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9382w9579w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9382w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9388w9587w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9388w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9394w9595w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9394w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9400w9603w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9400w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9406w9611w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9406w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9410w9619w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9410w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9304w9475w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9304w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9238w9627w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9238w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9243w9635w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9243w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9245w9643w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9245w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9247w9651w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9247w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9249w9659w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9249w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9251w9667w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9251w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9253w9675w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9253w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9255w9683w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9255w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9257w9691w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9257w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9259w9699w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9259w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9310w9483w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9310w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9261w9707w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9261w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9263w9715w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9263w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9316w9491w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9316w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9322w9499w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9322w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9328w9507w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9328w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9334w9515w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9334w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9340w9523w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9340w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9346w9531w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9346w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9352w9539w(0) <= wire_ccc_cordic_m_w_x_prenodeone_13_w_range9352w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range719w984w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range719w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range778w1066w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range778w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range784w1074w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range784w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range790w1082w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range790w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range796w1090w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range796w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range802w1098w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range802w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range808w1106w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range808w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range814w1114w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range814w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range820w1122w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range820w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range826w1130w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range826w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range832w1138w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range832w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range724w994w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range724w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range838w1146w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range838w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range844w1154w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range844w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range850w1162w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range850w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range856w1170w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range856w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range862w1178w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range862w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range868w1186w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range868w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range874w1194w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range874w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range880w1202w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range880w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range886w1210w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range886w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range892w1218w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range892w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range730w1002w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range730w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range896w1226w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range896w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range702w1234w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range702w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range736w1010w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range736w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range742w1018w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range742w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range748w1026w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range748w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range754w1034w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range754w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range760w1042w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range760w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range766w1050w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range766w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range772w1058w(0) <= wire_ccc_cordic_m_w_x_prenodeone_2_w_range772w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1524w1780w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1524w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1583w1862w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1583w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1589w1870w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1589w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1595w1878w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1595w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1601w1886w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1601w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1607w1894w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1607w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1613w1902w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1613w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1619w1910w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1619w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1625w1918w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1625w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1631w1926w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1631w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1637w1934w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1637w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1529w1790w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1529w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1643w1942w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1643w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1649w1950w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1649w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1655w1958w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1655w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1661w1966w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1661w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1667w1974w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1667w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1673w1982w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1673w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1679w1990w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1679w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1685w1998w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1685w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1691w2006w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1691w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1695w2014w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1695w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1535w1798w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1535w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1503w2022w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1503w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1508w2030w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1508w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1541w1806w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1541w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1547w1814w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1547w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1553w1822w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1553w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1559w1830w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1559w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1565w1838w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1565w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1571w1846w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1571w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1577w1854w(0) <= wire_ccc_cordic_m_w_x_prenodeone_3_w_range1577w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2324w2571w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2324w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2383w2653w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2383w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2389w2661w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2389w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2395w2669w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2395w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2401w2677w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2401w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2407w2685w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2407w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2413w2693w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2413w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2419w2701w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2419w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2425w2709w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2425w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2431w2717w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2431w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2437w2725w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2437w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2329w2581w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2329w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2443w2733w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2443w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2449w2741w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2449w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2455w2749w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2455w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2461w2757w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2461w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2467w2765w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2467w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2473w2773w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2473w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2479w2781w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2479w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2485w2789w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2485w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2489w2797w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2489w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2299w2805w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2299w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2335w2589w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2335w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2304w2813w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2304w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2306w2821w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2306w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2341w2597w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2341w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2347w2605w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2347w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2353w2613w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2353w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2359w2621w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2359w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2365w2629w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2365w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2371w2637w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2371w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2377w2645w(0) <= wire_ccc_cordic_m_w_x_prenodeone_4_w_range2377w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3119w3357w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3119w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3178w3439w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3178w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3184w3447w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3184w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3190w3455w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3190w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3196w3463w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3196w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3202w3471w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3202w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3208w3479w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3208w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3214w3487w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3214w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3220w3495w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3220w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3226w3503w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3226w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3232w3511w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3232w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3124w3367w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3124w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3238w3519w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3238w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3244w3527w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3244w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3250w3535w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3250w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3256w3543w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3256w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3262w3551w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3262w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3268w3559w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3268w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3274w3567w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3274w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3278w3575w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3278w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3090w3583w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3090w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3095w3591w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3095w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3130w3375w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3130w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3097w3599w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3097w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3099w3607w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3099w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3136w3383w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3136w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3142w3391w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3142w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3148w3399w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3148w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3154w3407w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3154w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3160w3415w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3160w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3166w3423w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3166w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3172w3431w(0) <= wire_ccc_cordic_m_w_x_prenodeone_5_w_range3172w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3909w4138w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3909w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3968w4220w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3968w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3974w4228w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3974w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3980w4236w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3980w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3986w4244w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3986w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3992w4252w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3992w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3998w4260w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3998w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4004w4268w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4004w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4010w4276w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4010w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4016w4284w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4016w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4022w4292w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4022w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3914w4148w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3914w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4028w4300w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4028w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4034w4308w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4034w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4040w4316w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4040w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4046w4324w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4046w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4052w4332w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4052w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4058w4340w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4058w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4062w4348w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range4062w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3876w4356w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3876w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3881w4364w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3881w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3883w4372w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3883w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3920w4156w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3920w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3885w4380w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3885w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3887w4388w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3887w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3926w4164w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3926w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3932w4172w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3932w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3938w4180w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3938w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3944w4188w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3944w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3950w4196w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3950w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3956w4204w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3956w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3962w4212w(0) <= wire_ccc_cordic_m_w_x_prenodeone_6_w_range3962w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4694w4914w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4694w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4753w4996w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4753w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4759w5004w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4759w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4765w5012w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4765w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4771w5020w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4771w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4777w5028w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4777w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4783w5036w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4783w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4789w5044w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4789w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4795w5052w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4795w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4801w5060w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4801w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4807w5068w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4807w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4699w4924w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4699w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4813w5076w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4813w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4819w5084w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4819w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4825w5092w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4825w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4831w5100w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4831w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4837w5108w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4837w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4841w5116w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4841w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4657w5124w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4657w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4662w5132w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4662w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4664w5140w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4664w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4666w5148w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4666w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4705w4932w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4705w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4668w5156w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4668w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4670w5164w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4670w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4711w4940w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4711w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4717w4948w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4717w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4723w4956w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4723w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4729w4964w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4729w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4735w4972w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4735w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4741w4980w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4741w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4747w4988w(0) <= wire_ccc_cordic_m_w_x_prenodeone_7_w_range4747w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5474w5685w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5474w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5533w5767w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5533w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5539w5775w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5539w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5545w5783w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5545w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5551w5791w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5551w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5557w5799w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5557w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5563w5807w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5563w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5569w5815w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5569w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5575w5823w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5575w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5581w5831w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5581w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5587w5839w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5587w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5479w5695w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5479w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5593w5847w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5593w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5599w5855w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5599w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5605w5863w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5605w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5611w5871w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5611w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5615w5879w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5615w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5433w5887w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5433w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5438w5895w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5438w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5440w5903w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5440w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5442w5911w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5442w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5444w5919w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5444w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5485w5703w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5485w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5446w5927w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5446w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5448w5935w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5448w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5491w5711w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5491w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5497w5719w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5497w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5503w5727w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5503w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5509w5735w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5509w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5515w5743w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5515w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5521w5751w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5521w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5527w5759w(0) <= wire_ccc_cordic_m_w_x_prenodeone_8_w_range5527w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6249w6451w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6249w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6308w6533w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6308w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6314w6541w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6314w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6320w6549w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6320w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6326w6557w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6326w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6332w6565w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6332w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6338w6573w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6338w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6344w6581w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6344w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6350w6589w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6350w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6356w6597w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6356w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6362w6605w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6362w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6254w6461w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6254w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6368w6613w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6368w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6374w6621w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6374w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6380w6629w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6380w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6384w6637w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6384w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6204w6645w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6204w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6209w6653w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6209w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6211w6661w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6211w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6213w6669w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6213w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6215w6677w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6215w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6217w6685w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6217w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6260w6469w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6260w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6219w6693w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6219w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6221w6701w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6221w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6266w6477w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6266w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6272w6485w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6272w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6278w6493w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6278w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6284w6501w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6284w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6290w6509w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6290w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6296w6517w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6296w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6302w6525w(0) <= wire_ccc_cordic_m_w_x_prenodeone_9_w_range6302w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7151w7210w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7151w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7180w7293w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7180w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7183w7301w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7183w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7186w7309w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7186w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7189w7317w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7189w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7192w7325w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7192w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7195w7333w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7195w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7198w7341w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7198w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7201w7349w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7201w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7204w7357w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7204w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7207w7365w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7207w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7153w7221w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7153w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range6991w7373w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range6991w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range6995w7381w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range6995w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range6997w7389w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range6997w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range6999w7397w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range6999w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7001w7405w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7001w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7003w7413w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7003w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7005w7421w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7005w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7007w7429w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7007w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7009w7437w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7009w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7011w7445w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7011w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7156w7229w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7156w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7013w7453w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7013w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7015w7461w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7015w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7159w7237w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7159w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7162w7245w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7162w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7165w7253w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7165w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7168w7261w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7168w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7171w7269w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7171w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7174w7277w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7174w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7177w7285w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7177w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7910w7966w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7910w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7939w8049w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7939w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7942w8057w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7942w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7945w8065w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7945w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7948w8073w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7948w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7951w8081w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7951w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7954w8089w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7954w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7957w8097w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7957w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7960w8105w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7960w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7963w8113w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7963w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7754w8121w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7754w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7912w7977w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7912w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7758w8129w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7758w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7760w8137w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7760w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7762w8145w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7762w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7764w8153w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7764w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7766w8161w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7766w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7768w8169w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7768w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7770w8177w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7770w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7772w8185w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7772w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7774w8193w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7774w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7776w8201w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7776w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7915w7985w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7915w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7778w8209w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7778w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7780w8217w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7780w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7918w7993w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7918w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7921w8001w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7921w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7924w8009w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7924w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7927w8017w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7927w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7930w8025w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7930w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7933w8033w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7933w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7936w8041w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7936w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8664w8717w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8664w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8693w8800w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8693w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8696w8808w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8696w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8699w8816w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8699w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8702w8824w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8702w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8705w8832w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8705w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8708w8840w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8708w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8711w8848w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8711w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8714w8856w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8714w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8512w8864w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8512w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8516w8872w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8516w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8666w8728w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8666w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8518w8880w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8518w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8520w8888w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8520w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8522w8896w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8522w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8524w8904w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8524w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8526w8912w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8526w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8528w8920w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8528w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8530w8928w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8530w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8532w8936w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8532w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8534w8944w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8534w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8536w8952w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8536w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8669w8736w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8669w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8538w8960w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8538w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8540w8968w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8540w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8672w8744w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8672w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8675w8752w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8675w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8678w8760w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8678w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8681w8768w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8681w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8684w8776w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8684w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8687w8784w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8687w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8690w8792w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8690w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9413w9463w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9413w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9442w9546w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9442w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9445w9554w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9445w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9448w9562w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9448w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9451w9570w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9451w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9454w9578w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9454w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9457w9586w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9457w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9460w9594w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9460w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9265w9602w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9265w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9269w9610w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9269w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9271w9618w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9271w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9415w9474w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9415w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9273w9626w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9273w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9275w9634w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9275w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9277w9642w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9277w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9279w9650w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9279w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9281w9658w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9281w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9283w9666w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9283w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9285w9674w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9285w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9287w9682w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9287w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9289w9690w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9289w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9291w9698w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9291w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9418w9482w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9418w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9293w9706w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9293w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9295w9714w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9295w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9421w9490w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9421w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9424w9498w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9424w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9427w9506w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9427w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9430w9514w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9430w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9433w9522w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9433w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9436w9530w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9436w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9439w9538w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9439w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range899w982w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range899w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range928w1065w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range928w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range931w1073w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range931w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range934w1081w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range934w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range937w1089w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range937w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range940w1097w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range940w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range943w1105w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range943w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range946w1113w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range946w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range949w1121w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range949w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range952w1129w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range952w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range955w1137w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range955w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range901w993w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range901w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range958w1145w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range958w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range961w1153w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range961w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range964w1161w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range964w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range967w1169w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range967w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range970w1177w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range970w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range973w1185w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range973w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range976w1193w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range976w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range979w1201w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range979w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range707w1209w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range707w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range711w1217w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range711w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range904w1001w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range904w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range713w1225w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range713w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range715w1233w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range715w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range907w1009w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range907w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range910w1017w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range910w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range913w1025w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range913w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range916w1033w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range916w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range919w1041w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range919w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range922w1049w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range922w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range925w1057w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_2_w_range925w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1698w1778w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1698w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1727w1861w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1727w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1730w1869w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1730w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1733w1877w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1733w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1736w1885w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1736w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1739w1893w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1739w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1742w1901w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1742w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1745w1909w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1745w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1748w1917w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1748w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1751w1925w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1751w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1754w1933w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1754w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1700w1789w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1700w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1757w1941w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1757w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1760w1949w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1760w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1763w1957w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1763w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1766w1965w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1766w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1769w1973w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1769w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1772w1981w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1772w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1775w1989w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1775w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1510w1997w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1510w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1514w2005w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1514w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1516w2013w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1516w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1703w1797w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1703w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1518w2021w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1518w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1520w2029w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1520w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1706w1805w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1706w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1709w1813w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1709w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1712w1821w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1712w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1715w1829w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1715w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1718w1837w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1718w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1721w1845w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1721w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1724w1853w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1724w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2492w2569w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2492w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2521w2652w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2521w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2524w2660w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2524w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2527w2668w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2527w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2530w2676w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2530w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2533w2684w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2533w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2536w2692w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2536w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2539w2700w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2539w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2542w2708w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2542w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2545w2716w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2545w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2548w2724w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2548w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2494w2580w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2494w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2551w2732w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2551w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2554w2740w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2554w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2557w2748w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2557w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2560w2756w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2560w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2563w2764w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2563w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2566w2772w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2566w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2308w2780w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2308w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2312w2788w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2312w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2314w2796w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2314w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2316w2804w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2316w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2497w2588w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2497w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2318w2812w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2318w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2320w2820w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2320w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2500w2596w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2500w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2503w2604w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2503w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2506w2612w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2506w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2509w2620w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2509w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2512w2628w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2512w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2515w2636w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2515w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2518w2644w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2518w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3281w3355w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3281w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3310w3438w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3310w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3313w3446w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3313w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3316w3454w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3316w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3319w3462w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3319w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3322w3470w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3322w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3325w3478w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3325w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3328w3486w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3328w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3331w3494w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3331w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3334w3502w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3334w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3337w3510w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3337w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3283w3366w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3283w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3340w3518w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3340w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3343w3526w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3343w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3346w3534w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3346w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3349w3542w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3349w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3352w3550w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3352w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3101w3558w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3101w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3105w3566w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3105w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3107w3574w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3107w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3109w3582w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3109w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3111w3590w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3111w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3286w3374w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3286w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3113w3598w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3113w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3115w3606w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3115w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3289w3382w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3289w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3292w3390w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3292w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3295w3398w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3295w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3298w3406w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3298w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3301w3414w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3301w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3304w3422w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3304w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3307w3430w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3307w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4065w4136w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4065w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4094w4219w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4094w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4097w4227w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4097w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4100w4235w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4100w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4103w4243w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4103w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4106w4251w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4106w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4109w4259w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4109w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4112w4267w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4112w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4115w4275w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4115w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4118w4283w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4118w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4121w4291w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4121w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4067w4147w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4067w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4124w4299w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4124w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4127w4307w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4127w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4130w4315w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4130w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4133w4323w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4133w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3889w4331w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3889w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3893w4339w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3893w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3895w4347w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3895w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3897w4355w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3897w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3899w4363w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3899w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3901w4371w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3901w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4070w4155w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4070w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3903w4379w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3903w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3905w4387w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3905w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4073w4163w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4073w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4076w4171w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4076w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4079w4179w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4079w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4082w4187w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4082w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4085w4195w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4085w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4088w4203w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4088w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4091w4211w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4091w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4844w4912w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4844w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4873w4995w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4873w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4876w5003w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4876w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4879w5011w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4879w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4882w5019w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4882w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4885w5027w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4885w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4888w5035w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4888w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4891w5043w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4891w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4894w5051w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4894w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4897w5059w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4897w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4900w5067w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4900w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4846w4923w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4846w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4903w5075w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4903w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4906w5083w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4906w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4909w5091w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4909w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4672w5099w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4672w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4676w5107w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4676w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4678w5115w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4678w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4680w5123w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4680w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4682w5131w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4682w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4684w5139w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4684w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4686w5147w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4686w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4849w4931w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4849w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4688w5155w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4688w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4690w5163w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4690w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4852w4939w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4852w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4855w4947w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4855w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4858w4955w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4858w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4861w4963w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4861w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4864w4971w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4864w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4867w4979w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4867w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4870w4987w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4870w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5618w5683w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5618w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5647w5766w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5647w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5650w5774w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5650w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5653w5782w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5653w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5656w5790w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5656w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5659w5798w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5659w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5662w5806w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5662w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5665w5814w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5665w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5668w5822w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5668w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5671w5830w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5671w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5674w5838w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5674w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5620w5694w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5620w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5677w5846w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5677w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5680w5854w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5680w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5450w5862w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5450w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5454w5870w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5454w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5456w5878w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5456w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5458w5886w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5458w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5460w5894w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5460w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5462w5902w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5462w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5464w5910w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5464w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5466w5918w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5466w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5623w5702w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5623w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5468w5926w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5468w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5470w5934w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5470w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5626w5710w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5626w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5629w5718w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5629w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5632w5726w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5632w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5635w5734w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5635w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5638w5742w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5638w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5641w5750w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5641w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5644w5758w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5644w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6387w6449w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6387w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6416w6532w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6416w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6419w6540w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6419w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6422w6548w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6422w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6425w6556w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6425w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6428w6564w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6428w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6431w6572w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6431w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6434w6580w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6434w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6437w6588w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6437w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6440w6596w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6440w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6443w6604w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6443w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6389w6460w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6389w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6446w6612w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6446w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6223w6620w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6223w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6227w6628w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6227w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6229w6636w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6229w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6231w6644w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6231w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6233w6652w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6233w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6235w6660w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6235w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6237w6668w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6237w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6239w6676w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6239w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6241w6684w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6241w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6392w6468w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6392w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6243w6692w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6243w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6245w6700w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6245w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6395w6476w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6395w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6398w6484w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6398w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6401w6492w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6401w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6404w6500w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6404w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6407w6508w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6407w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6410w6516w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6410w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6413w6524w(0) <= wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6413w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7021w7217w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7021w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7080w7298w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7080w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7086w7306w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7086w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7092w7314w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7092w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7098w7322w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7098w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7104w7330w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7104w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7110w7338w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7110w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7116w7346w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7116w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7122w7354w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7122w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7128w7362w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7128w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7134w7370w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7134w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7026w7226w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7026w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7140w7378w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7140w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7146w7386w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7146w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7149w7394w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7149w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6973w7402w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range6973w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6976w7410w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range6976w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6978w7418w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range6978w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6980w7426w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range6980w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6982w7434w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range6982w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6984w7442w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range6984w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6986w7450w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range6986w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7032w7234w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7032w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6988w7458w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range6988w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6990w7466w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range6990w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7038w7242w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7038w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7044w7250w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7044w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7050w7258w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7050w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7056w7266w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7056w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7062w7274w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7062w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7068w7282w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7068w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7074w7290w(0) <= wire_ccc_cordic_m_w_y_prenodeone_10_w_range7074w(0) AND wire_indexbitff_w_lg_w_q_range474w7211w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7786w7973w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7786w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7845w8054w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7845w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7851w8062w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7851w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7857w8070w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7857w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7863w8078w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7863w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7869w8086w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7869w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7875w8094w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7875w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7881w8102w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7881w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7887w8110w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7887w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7893w8118w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7893w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7899w8126w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7899w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7791w7982w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7791w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7905w8134w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7905w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7908w8142w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7908w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7734w8150w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7734w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7737w8158w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7737w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7739w8166w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7739w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7741w8174w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7741w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7743w8182w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7743w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7745w8190w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7745w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7747w8198w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7747w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7749w8206w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7749w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7797w7990w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7797w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7751w8214w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7751w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7753w8222w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7753w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7803w7998w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7803w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7809w8006w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7809w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7815w8014w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7815w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7821w8022w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7821w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7827w8030w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7827w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7833w8038w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7833w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7839w8046w(0) <= wire_ccc_cordic_m_w_y_prenodeone_11_w_range7839w(0) AND wire_indexbitff_w_lg_w_q_range477w7967w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8546w8724w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8546w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8605w8805w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8605w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8611w8813w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8611w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8617w8821w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8617w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8623w8829w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8623w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8629w8837w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8629w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8635w8845w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8635w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8641w8853w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8641w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8647w8861w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8647w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8653w8869w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8653w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8659w8877w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8659w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8551w8733w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8551w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8662w8885w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8662w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8490w8893w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8490w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8493w8901w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8493w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8495w8909w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8495w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8497w8917w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8497w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8499w8925w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8499w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8501w8933w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8501w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8503w8941w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8503w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8505w8949w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8505w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8507w8957w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8507w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8557w8741w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8557w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8509w8965w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8509w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8511w8973w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8511w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8563w8749w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8563w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8569w8757w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8569w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8575w8765w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8575w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8581w8773w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8581w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8587w8781w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8587w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8593w8789w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8593w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8599w8797w(0) <= wire_ccc_cordic_m_w_y_prenodeone_12_w_range8599w(0) AND wire_indexbitff_w_lg_w_q_range480w8718w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9301w9470w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9301w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9360w9551w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9360w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9366w9559w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9366w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9372w9567w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9372w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9378w9575w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9378w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9384w9583w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9384w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9390w9591w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9390w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9396w9599w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9396w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9402w9607w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9402w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9408w9615w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9408w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9411w9623w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9411w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9306w9479w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9306w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9241w9631w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9241w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9244w9639w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9244w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9246w9647w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9246w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9248w9655w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9248w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9250w9663w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9250w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9252w9671w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9252w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9254w9679w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9254w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9256w9687w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9256w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9258w9695w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9258w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9260w9703w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9260w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9312w9487w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9312w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9262w9711w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9262w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9264w9719w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9264w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9318w9495w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9318w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9324w9503w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9324w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9330w9511w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9330w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9336w9519w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9336w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9342w9527w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9342w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9348w9535w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9348w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9354w9543w(0) <= wire_ccc_cordic_m_w_y_prenodeone_13_w_range9354w(0) AND wire_indexbitff_w_lg_w_q_range483w9464w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range721w989w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range721w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range780w1070w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range780w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range786w1078w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range786w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range792w1086w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range792w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range798w1094w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range798w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range804w1102w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range804w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range810w1110w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range810w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range816w1118w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range816w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range822w1126w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range822w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range828w1134w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range828w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range834w1142w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range834w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range726w998w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range726w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range840w1150w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range840w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range846w1158w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range846w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range852w1166w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range852w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range858w1174w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range858w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range864w1182w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range864w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range870w1190w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range870w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range876w1198w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range876w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range882w1206w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range882w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range888w1214w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range888w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range894w1222w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range894w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range732w1006w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range732w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range897w1230w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range897w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range705w1238w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range705w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range738w1014w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range738w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range744w1022w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range744w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range750w1030w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range750w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range756w1038w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range756w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range762w1046w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range762w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range768w1054w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range768w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range774w1062w(0) <= wire_ccc_cordic_m_w_y_prenodeone_2_w_range774w(0) AND wire_indexbitff_w_lg_w_q_range450w983w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1526w1785w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1526w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1585w1866w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1585w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1591w1874w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1591w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1597w1882w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1597w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1603w1890w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1603w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1609w1898w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1609w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1615w1906w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1615w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1621w1914w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1621w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1627w1922w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1627w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1633w1930w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1633w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1639w1938w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1639w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1531w1794w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1531w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1645w1946w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1645w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1651w1954w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1651w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1657w1962w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1657w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1663w1970w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1663w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1669w1978w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1669w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1675w1986w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1675w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1681w1994w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1681w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1687w2002w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1687w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1693w2010w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1693w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1696w2018w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1696w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1537w1802w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1537w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1506w2026w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1506w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1509w2034w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1509w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1543w1810w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1543w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1549w1818w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1549w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1555w1826w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1555w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1561w1834w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1561w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1567w1842w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1567w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1573w1850w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1573w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1579w1858w(0) <= wire_ccc_cordic_m_w_y_prenodeone_3_w_range1579w(0) AND wire_indexbitff_w_lg_w_q_range453w1779w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2326w2576w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2326w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2385w2657w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2385w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2391w2665w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2391w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2397w2673w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2397w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2403w2681w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2403w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2409w2689w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2409w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2415w2697w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2415w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2421w2705w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2421w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2427w2713w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2427w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2433w2721w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2433w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2439w2729w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2439w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2331w2585w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2331w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2445w2737w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2445w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2451w2745w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2451w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2457w2753w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2457w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2463w2761w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2463w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2469w2769w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2469w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2475w2777w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2475w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2481w2785w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2481w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2487w2793w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2487w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2490w2801w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2490w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2302w2809w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2302w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2337w2593w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2337w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2305w2817w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2305w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2307w2825w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2307w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2343w2601w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2343w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2349w2609w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2349w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2355w2617w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2355w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2361w2625w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2361w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2367w2633w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2367w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2373w2641w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2373w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2379w2649w(0) <= wire_ccc_cordic_m_w_y_prenodeone_4_w_range2379w(0) AND wire_indexbitff_w_lg_w_q_range456w2570w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3121w3362w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3121w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3180w3443w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3180w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3186w3451w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3186w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3192w3459w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3192w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3198w3467w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3198w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3204w3475w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3204w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3210w3483w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3210w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3216w3491w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3216w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3222w3499w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3222w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3228w3507w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3228w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3234w3515w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3234w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3126w3371w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3126w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3240w3523w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3240w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3246w3531w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3246w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3252w3539w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3252w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3258w3547w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3258w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3264w3555w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3264w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3270w3563w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3270w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3276w3571w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3276w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3279w3579w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3279w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3093w3587w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3093w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3096w3595w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3096w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3132w3379w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3132w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3098w3603w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3098w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3100w3611w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3100w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3138w3387w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3138w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3144w3395w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3144w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3150w3403w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3150w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3156w3411w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3156w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3162w3419w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3162w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3168w3427w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3168w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3174w3435w(0) <= wire_ccc_cordic_m_w_y_prenodeone_5_w_range3174w(0) AND wire_indexbitff_w_lg_w_q_range459w3356w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3911w4143w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3911w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3970w4224w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3970w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3976w4232w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3976w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3982w4240w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3982w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3988w4248w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3988w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3994w4256w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3994w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4000w4264w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4000w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4006w4272w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4006w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4012w4280w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4012w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4018w4288w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4018w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4024w4296w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4024w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3916w4152w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3916w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4030w4304w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4030w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4036w4312w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4036w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4042w4320w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4042w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4048w4328w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4048w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4054w4336w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4054w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4060w4344w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4060w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4063w4352w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range4063w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3879w4360w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3879w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3882w4368w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3882w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3884w4376w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3884w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3922w4160w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3922w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3886w4384w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3886w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3888w4392w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3888w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3928w4168w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3928w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3934w4176w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3934w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3940w4184w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3940w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3946w4192w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3946w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3952w4200w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3952w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3958w4208w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3958w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3964w4216w(0) <= wire_ccc_cordic_m_w_y_prenodeone_6_w_range3964w(0) AND wire_indexbitff_w_lg_w_q_range462w4137w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4696w4919w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4696w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4755w5000w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4755w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4761w5008w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4761w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4767w5016w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4767w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4773w5024w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4773w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4779w5032w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4779w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4785w5040w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4785w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4791w5048w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4791w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4797w5056w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4797w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4803w5064w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4803w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4809w5072w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4809w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4701w4928w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4701w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4815w5080w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4815w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4821w5088w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4821w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4827w5096w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4827w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4833w5104w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4833w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4839w5112w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4839w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4842w5120w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4842w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4660w5128w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4660w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4663w5136w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4663w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4665w5144w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4665w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4667w5152w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4667w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4707w4936w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4707w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4669w5160w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4669w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4671w5168w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4671w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4713w4944w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4713w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4719w4952w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4719w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4725w4960w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4725w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4731w4968w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4731w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4737w4976w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4737w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4743w4984w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4743w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4749w4992w(0) <= wire_ccc_cordic_m_w_y_prenodeone_7_w_range4749w(0) AND wire_indexbitff_w_lg_w_q_range465w4913w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5476w5690w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5476w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5535w5771w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5535w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5541w5779w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5541w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5547w5787w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5547w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5553w5795w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5553w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5559w5803w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5559w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5565w5811w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5565w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5571w5819w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5571w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5577w5827w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5577w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5583w5835w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5583w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5589w5843w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5589w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5481w5699w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5481w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5595w5851w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5595w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5601w5859w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5601w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5607w5867w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5607w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5613w5875w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5613w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5616w5883w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5616w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5436w5891w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5436w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5439w5899w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5439w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5441w5907w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5441w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5443w5915w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5443w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5445w5923w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5445w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5487w5707w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5487w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5447w5931w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5447w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5449w5939w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5449w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5493w5715w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5493w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5499w5723w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5499w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5505w5731w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5505w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5511w5739w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5511w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5517w5747w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5517w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5523w5755w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5523w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5529w5763w(0) <= wire_ccc_cordic_m_w_y_prenodeone_8_w_range5529w(0) AND wire_indexbitff_w_lg_w_q_range468w5684w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6251w6456w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6251w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6310w6537w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6310w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6316w6545w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6316w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6322w6553w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6322w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6328w6561w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6328w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6334w6569w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6334w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6340w6577w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6340w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6346w6585w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6346w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6352w6593w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6352w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6358w6601w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6358w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6364w6609w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6364w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6256w6465w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6256w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6370w6617w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6370w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6376w6625w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6376w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6382w6633w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6382w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6385w6641w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6385w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6207w6649w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6207w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6210w6657w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6210w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6212w6665w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6212w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6214w6673w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6214w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6216w6681w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6216w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6218w6689w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6218w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6262w6473w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6262w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6220w6697w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6220w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6222w6705w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6222w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6268w6481w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6268w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6274w6489w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6274w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6280w6497w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6280w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6286w6505w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6286w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6292w6513w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6292w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6298w6521w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6298w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6304w6529w(0) <= wire_ccc_cordic_m_w_y_prenodeone_9_w_range6304w(0) AND wire_indexbitff_w_lg_w_q_range471w6450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7152w7216w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7152w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7181w7297w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7181w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7184w7305w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7184w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7187w7313w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7187w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7190w7321w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7190w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7193w7329w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7193w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7196w7337w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7196w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7199w7345w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7199w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7202w7353w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7202w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7205w7361w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7205w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7208w7369w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7208w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7154w7225w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7154w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range6993w7377w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range6993w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range6996w7385w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range6996w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range6998w7393w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range6998w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7000w7401w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7000w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7002w7409w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7002w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7004w7417w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7004w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7006w7425w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7006w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7008w7433w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7008w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7010w7441w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7010w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7012w7449w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7012w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7157w7233w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7157w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7014w7457w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7014w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7016w7465w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7016w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7160w7241w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7160w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7163w7249w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7163w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7166w7257w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7166w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7169w7265w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7169w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7172w7273w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7172w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7175w7281w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7175w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7178w7289w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7178w(0) AND wire_indexbitff_w_q_range474w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7911w7972w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7911w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7940w8053w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7940w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7943w8061w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7943w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7946w8069w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7946w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7949w8077w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7949w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7952w8085w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7952w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7955w8093w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7955w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7958w8101w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7958w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7961w8109w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7961w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7964w8117w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7964w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7756w8125w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7756w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7913w7981w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7913w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7759w8133w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7759w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7761w8141w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7761w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7763w8149w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7763w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7765w8157w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7765w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7767w8165w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7767w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7769w8173w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7769w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7771w8181w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7771w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7773w8189w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7773w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7775w8197w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7775w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7777w8205w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7777w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7916w7989w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7916w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7779w8213w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7779w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7781w8221w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7781w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7919w7997w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7919w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7922w8005w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7922w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7925w8013w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7925w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7928w8021w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7928w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7931w8029w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7931w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7934w8037w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7934w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7937w8045w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7937w(0) AND wire_indexbitff_w_q_range477w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8665w8723w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8665w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8694w8804w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8694w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8697w8812w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8697w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8700w8820w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8700w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8703w8828w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8703w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8706w8836w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8706w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8709w8844w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8709w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8712w8852w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8712w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8715w8860w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8715w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8514w8868w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8514w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8517w8876w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8517w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8667w8732w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8667w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8519w8884w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8519w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8521w8892w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8521w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8523w8900w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8523w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8525w8908w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8525w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8527w8916w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8527w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8529w8924w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8529w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8531w8932w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8531w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8533w8940w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8533w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8535w8948w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8535w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8537w8956w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8537w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8670w8740w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8670w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8539w8964w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8539w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8541w8972w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8541w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8673w8748w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8673w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8676w8756w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8676w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8679w8764w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8679w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8682w8772w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8682w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8685w8780w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8685w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8688w8788w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8688w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8691w8796w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8691w(0) AND wire_indexbitff_w_q_range480w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9414w9469w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9414w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9443w9550w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9443w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9446w9558w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9446w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9449w9566w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9449w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9452w9574w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9452w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9455w9582w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9455w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9458w9590w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9458w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9461w9598w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9461w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9267w9606w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9267w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9270w9614w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9270w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9272w9622w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9272w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9416w9478w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9416w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9274w9630w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9274w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9276w9638w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9276w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9278w9646w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9278w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9280w9654w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9280w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9282w9662w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9282w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9284w9670w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9284w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9286w9678w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9286w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9288w9686w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9288w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9290w9694w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9290w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9292w9702w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9292w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9419w9486w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9419w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9294w9710w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9294w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9296w9718w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9296w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9422w9494w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9422w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9425w9502w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9425w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9428w9510w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9428w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9431w9518w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9431w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9434w9526w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9434w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9437w9534w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9437w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9440w9542w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9440w(0) AND wire_indexbitff_w_q_range483w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range900w988w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range900w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range929w1069w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range929w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range932w1077w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range932w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range935w1085w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range935w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range938w1093w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range938w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range941w1101w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range941w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range944w1109w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range944w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range947w1117w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range947w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range950w1125w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range950w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range953w1133w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range953w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range956w1141w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range956w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range902w997w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range902w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range959w1149w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range959w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range962w1157w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range962w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range965w1165w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range965w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range968w1173w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range968w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range971w1181w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range971w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range974w1189w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range974w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range977w1197w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range977w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range980w1205w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range980w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range709w1213w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range709w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range712w1221w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range712w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range905w1005w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range905w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range714w1229w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range714w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range716w1237w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range716w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range908w1013w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range908w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range911w1021w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range911w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range914w1029w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range914w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range917w1037w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range917w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range920w1045w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range920w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range923w1053w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range923w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range926w1061w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_2_w_range926w(0) AND wire_indexbitff_w_q_range450w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1699w1784w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1699w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1728w1865w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1728w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1731w1873w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1731w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1734w1881w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1734w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1737w1889w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1737w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1740w1897w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1740w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1743w1905w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1743w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1746w1913w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1746w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1749w1921w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1749w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1752w1929w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1752w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1755w1937w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1755w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1701w1793w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1701w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1758w1945w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1758w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1761w1953w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1761w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1764w1961w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1764w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1767w1969w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1767w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1770w1977w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1770w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1773w1985w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1773w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1776w1993w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1776w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1512w2001w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1512w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1515w2009w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1515w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1517w2017w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1517w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1704w1801w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1704w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1519w2025w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1519w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1521w2033w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1521w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1707w1809w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1707w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1710w1817w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1710w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1713w1825w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1713w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1716w1833w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1716w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1719w1841w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1719w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1722w1849w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1722w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1725w1857w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1725w(0) AND wire_indexbitff_w_q_range453w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2493w2575w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2493w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2522w2656w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2522w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2525w2664w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2525w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2528w2672w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2528w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2531w2680w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2531w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2534w2688w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2534w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2537w2696w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2537w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2540w2704w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2540w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2543w2712w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2543w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2546w2720w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2546w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2549w2728w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2549w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2495w2584w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2495w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2552w2736w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2552w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2555w2744w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2555w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2558w2752w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2558w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2561w2760w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2561w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2564w2768w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2564w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2567w2776w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2567w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2310w2784w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2310w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2313w2792w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2313w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2315w2800w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2315w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2317w2808w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2317w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2498w2592w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2498w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2319w2816w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2319w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2321w2824w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2321w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2501w2600w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2501w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2504w2608w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2504w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2507w2616w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2507w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2510w2624w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2510w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2513w2632w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2513w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2516w2640w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2516w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2519w2648w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2519w(0) AND wire_indexbitff_w_q_range456w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3282w3361w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3282w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3311w3442w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3311w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3314w3450w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3314w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3317w3458w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3317w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3320w3466w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3320w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3323w3474w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3323w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3326w3482w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3326w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3329w3490w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3329w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3332w3498w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3332w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3335w3506w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3335w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3338w3514w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3338w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3284w3370w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3284w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3341w3522w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3341w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3344w3530w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3344w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3347w3538w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3347w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3350w3546w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3350w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3353w3554w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3353w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3103w3562w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3103w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3106w3570w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3106w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3108w3578w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3108w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3110w3586w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3110w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3112w3594w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3112w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3287w3378w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3287w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3114w3602w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3114w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3116w3610w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3116w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3290w3386w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3290w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3293w3394w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3293w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3296w3402w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3296w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3299w3410w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3299w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3302w3418w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3302w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3305w3426w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3305w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3308w3434w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3308w(0) AND wire_indexbitff_w_q_range459w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4066w4142w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4066w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4095w4223w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4095w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4098w4231w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4098w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4101w4239w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4101w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4104w4247w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4104w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4107w4255w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4107w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4110w4263w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4110w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4113w4271w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4113w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4116w4279w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4116w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4119w4287w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4119w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4122w4295w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4122w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4068w4151w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4068w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4125w4303w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4125w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4128w4311w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4128w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4131w4319w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4131w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4134w4327w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4134w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3891w4335w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3891w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3894w4343w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3894w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3896w4351w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3896w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3898w4359w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3898w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3900w4367w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3900w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3902w4375w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3902w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4071w4159w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4071w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3904w4383w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3904w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3906w4391w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3906w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4074w4167w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4074w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4077w4175w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4077w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4080w4183w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4080w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4083w4191w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4083w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4086w4199w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4086w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4089w4207w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4089w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4092w4215w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4092w(0) AND wire_indexbitff_w_q_range462w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4845w4918w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4845w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4874w4999w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4874w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4877w5007w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4877w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4880w5015w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4880w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4883w5023w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4883w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4886w5031w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4886w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4889w5039w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4889w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4892w5047w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4892w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4895w5055w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4895w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4898w5063w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4898w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4901w5071w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4901w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4847w4927w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4847w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4904w5079w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4904w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4907w5087w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4907w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4910w5095w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4910w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4674w5103w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4674w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4677w5111w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4677w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4679w5119w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4679w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4681w5127w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4681w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4683w5135w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4683w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4685w5143w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4685w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4687w5151w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4687w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4850w4935w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4850w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4689w5159w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4689w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4691w5167w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4691w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4853w4943w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4853w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4856w4951w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4856w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4859w4959w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4859w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4862w4967w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4862w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4865w4975w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4865w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4868w4983w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4868w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4871w4991w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4871w(0) AND wire_indexbitff_w_q_range465w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5619w5689w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5619w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5648w5770w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5648w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5651w5778w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5651w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5654w5786w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5654w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5657w5794w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5657w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5660w5802w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5660w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5663w5810w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5663w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5666w5818w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5666w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5669w5826w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5669w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5672w5834w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5672w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5675w5842w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5675w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5621w5698w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5621w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5678w5850w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5678w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5681w5858w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5681w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5452w5866w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5452w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5455w5874w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5455w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5457w5882w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5457w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5459w5890w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5459w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5461w5898w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5461w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5463w5906w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5463w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5465w5914w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5465w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5467w5922w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5467w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5624w5706w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5624w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5469w5930w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5469w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5471w5938w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5471w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5627w5714w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5627w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5630w5722w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5630w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5633w5730w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5633w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5636w5738w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5636w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5639w5746w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5639w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5642w5754w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5642w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5645w5762w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5645w(0) AND wire_indexbitff_w_q_range468w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6388w6455w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6388w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6417w6536w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6417w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6420w6544w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6420w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6423w6552w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6423w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6426w6560w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6426w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6429w6568w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6429w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6432w6576w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6432w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6435w6584w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6435w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6438w6592w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6438w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6441w6600w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6441w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6444w6608w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6444w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6390w6464w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6390w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6447w6616w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6447w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6225w6624w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6225w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6228w6632w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6228w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6230w6640w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6230w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6232w6648w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6232w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6234w6656w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6234w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6236w6664w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6236w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6238w6672w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6238w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6240w6680w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6240w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6242w6688w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6242w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6393w6472w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6393w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6244w6696w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6244w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6246w6704w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6246w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6396w6480w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6396w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6399w6488w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6399w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6402w6496w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6402w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6405w6504w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6405w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6408w6512w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6408w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6411w6520w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6411w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6414w6528w(0) <= wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6414w(0) AND wire_indexbitff_w_q_range471w(0);
	wire_ccc_cordic_m_w_lg_indexbit291w(0) <= NOT indexbit;
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8232w8233w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8232w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8313w8314w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8313w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8321w8322w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8321w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8329w8330w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8329w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8337w8338w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8337w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8345w8346w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8345w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8353w8354w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8353w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8361w8362w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8361w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8369w8370w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8369w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8377w8378w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8377w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8385w8386w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8385w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8241w8242w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8241w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8393w8394w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8393w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8401w8402w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8401w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8409w8410w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8409w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8417w8418w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8417w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8425w8426w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8425w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8433w8434w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8433w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8441w8442w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8441w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8449w8450w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8449w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8457w8458w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8457w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8465w8466w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8465w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8249w8250w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8249w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8473w8474w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8473w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8481w8482w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8481w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8257w8258w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8257w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8265w8266w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8265w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8273w8274w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8273w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8281w8282w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8281w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8289w8290w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8289w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8297w8298w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8297w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8305w8306w(0) <= NOT wire_ccc_cordic_m_w_atannode_10_w_range8305w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range8983w8984w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range8983w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9064w9065w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9064w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9072w9073w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9072w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9080w9081w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9080w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9088w9089w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9088w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9096w9097w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9096w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9104w9105w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9104w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9112w9113w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9112w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9120w9121w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9120w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9128w9129w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9128w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9136w9137w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9136w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range8992w8993w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range8992w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9144w9145w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9144w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9152w9153w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9152w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9160w9161w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9160w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9168w9169w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9168w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9176w9177w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9176w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9184w9185w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9184w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9192w9193w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9192w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9200w9201w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9200w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9208w9209w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9208w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9216w9217w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9216w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9000w9001w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9000w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9224w9225w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9224w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9232w9233w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9232w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9008w9009w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9008w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9016w9017w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9016w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9024w9025w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9024w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9032w9033w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9032w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9040w9041w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9040w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9048w9049w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9048w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9056w9057w(0) <= NOT wire_ccc_cordic_m_w_atannode_11_w_range9056w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9729w9730w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9729w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9810w9811w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9810w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9818w9819w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9818w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9826w9827w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9826w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9834w9835w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9834w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9842w9843w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9842w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9850w9851w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9850w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9858w9859w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9858w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9866w9867w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9866w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9874w9875w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9874w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9882w9883w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9882w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9738w9739w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9738w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9890w9891w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9890w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9898w9899w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9898w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9906w9907w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9906w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9914w9915w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9914w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9922w9923w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9922w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9930w9931w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9930w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9938w9939w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9938w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9946w9947w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9946w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9954w9955w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9954w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9962w9963w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9962w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9746w9747w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9746w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9970w9971w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9970w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9978w9979w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9978w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9754w9755w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9754w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9762w9763w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9762w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9770w9771w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9770w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9778w9779w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9778w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9786w9787w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9786w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9794w9795w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9794w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9802w9803w(0) <= NOT wire_ccc_cordic_m_w_atannode_12_w_range9802w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1248w1249w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1248w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1329w1330w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1329w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1337w1338w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1337w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1345w1346w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1345w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1353w1354w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1353w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1361w1362w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1361w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1369w1370w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1369w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1377w1378w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1377w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1385w1386w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1385w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1393w1394w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1393w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1401w1402w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1401w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1257w1258w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1257w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1409w1410w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1409w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1417w1418w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1417w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1425w1426w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1425w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1433w1434w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1433w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1441w1442w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1441w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1449w1450w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1449w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1457w1458w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1457w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1465w1466w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1465w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1473w1474w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1473w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1481w1482w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1481w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1265w1266w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1265w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1489w1490w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1489w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1497w1498w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1497w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1273w1274w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1273w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1281w1282w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1281w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1289w1290w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1289w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1297w1298w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1297w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1305w1306w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1305w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1313w1314w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1313w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1321w1322w(0) <= NOT wire_ccc_cordic_m_w_atannode_1_w_range1321w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2044w2045w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2044w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2125w2126w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2125w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2133w2134w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2133w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2141w2142w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2141w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2149w2150w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2149w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2157w2158w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2157w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2165w2166w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2165w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2173w2174w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2173w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2181w2182w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2181w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2189w2190w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2189w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2197w2198w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2197w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2053w2054w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2053w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2205w2206w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2205w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2213w2214w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2213w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2221w2222w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2221w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2229w2230w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2229w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2237w2238w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2237w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2245w2246w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2245w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2253w2254w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2253w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2261w2262w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2261w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2269w2270w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2269w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2277w2278w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2277w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2061w2062w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2061w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2285w2286w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2285w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2293w2294w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2293w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2069w2070w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2069w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2077w2078w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2077w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2085w2086w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2085w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2093w2094w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2093w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2101w2102w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2101w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2109w2110w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2109w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2117w2118w(0) <= NOT wire_ccc_cordic_m_w_atannode_2_w_range2117w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2835w2836w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2835w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2916w2917w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2916w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2924w2925w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2924w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2932w2933w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2932w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2940w2941w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2940w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2948w2949w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2948w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2956w2957w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2956w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2964w2965w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2964w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2972w2973w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2972w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2980w2981w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2980w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2988w2989w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2988w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2844w2845w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2844w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2996w2997w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2996w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3004w3005w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3004w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3012w3013w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3012w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3020w3021w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3020w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3028w3029w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3028w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3036w3037w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3036w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3044w3045w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3044w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3052w3053w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3052w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3060w3061w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3060w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3068w3069w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3068w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2852w2853w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2852w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3076w3077w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3076w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3084w3085w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range3084w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2860w2861w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2860w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2868w2869w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2868w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2876w2877w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2876w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2884w2885w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2884w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2892w2893w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2892w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2900w2901w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2900w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2908w2909w(0) <= NOT wire_ccc_cordic_m_w_atannode_3_w_range2908w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3621w3622w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3621w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3702w3703w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3702w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3710w3711w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3710w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3718w3719w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3718w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3726w3727w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3726w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3734w3735w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3734w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3742w3743w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3742w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3750w3751w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3750w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3758w3759w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3758w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3766w3767w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3766w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3774w3775w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3774w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3630w3631w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3630w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3782w3783w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3782w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3790w3791w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3790w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3798w3799w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3798w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3806w3807w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3806w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3814w3815w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3814w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3822w3823w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3822w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3830w3831w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3830w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3838w3839w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3838w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3846w3847w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3846w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3854w3855w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3854w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3638w3639w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3638w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3862w3863w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3862w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3870w3871w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3870w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3646w3647w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3646w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3654w3655w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3654w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3662w3663w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3662w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3670w3671w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3670w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3678w3679w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3678w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3686w3687w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3686w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3694w3695w(0) <= NOT wire_ccc_cordic_m_w_atannode_4_w_range3694w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4402w4403w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4402w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4483w4484w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4483w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4491w4492w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4491w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4499w4500w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4499w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4507w4508w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4507w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4515w4516w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4515w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4523w4524w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4523w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4531w4532w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4531w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4539w4540w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4539w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4547w4548w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4547w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4555w4556w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4555w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4411w4412w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4411w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4563w4564w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4563w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4571w4572w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4571w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4579w4580w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4579w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4587w4588w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4587w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4595w4596w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4595w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4603w4604w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4603w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4611w4612w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4611w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4619w4620w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4619w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4627w4628w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4627w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4635w4636w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4635w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4419w4420w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4419w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4643w4644w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4643w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4651w4652w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4651w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4427w4428w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4427w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4435w4436w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4435w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4443w4444w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4443w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4451w4452w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4451w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4459w4460w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4459w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4467w4468w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4467w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4475w4476w(0) <= NOT wire_ccc_cordic_m_w_atannode_5_w_range4475w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5178w5179w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5178w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5259w5260w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5259w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5267w5268w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5267w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5275w5276w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5275w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5283w5284w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5283w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5291w5292w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5291w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5299w5300w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5299w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5307w5308w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5307w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5315w5316w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5315w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5323w5324w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5323w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5331w5332w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5331w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5187w5188w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5187w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5339w5340w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5339w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5347w5348w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5347w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5355w5356w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5355w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5363w5364w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5363w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5371w5372w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5371w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5379w5380w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5379w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5387w5388w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5387w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5395w5396w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5395w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5403w5404w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5403w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5411w5412w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5411w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5195w5196w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5195w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5419w5420w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5419w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5427w5428w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5427w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5203w5204w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5203w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5211w5212w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5211w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5219w5220w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5219w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5227w5228w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5227w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5235w5236w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5235w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5243w5244w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5243w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5251w5252w(0) <= NOT wire_ccc_cordic_m_w_atannode_6_w_range5251w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5949w5950w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range5949w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6030w6031w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6030w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6038w6039w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6038w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6046w6047w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6046w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6054w6055w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6054w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6062w6063w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6062w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6070w6071w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6070w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6078w6079w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6078w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6086w6087w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6086w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6094w6095w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6094w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6102w6103w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6102w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5958w5959w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range5958w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6110w6111w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6110w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6118w6119w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6118w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6126w6127w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6126w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6134w6135w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6134w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6142w6143w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6142w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6150w6151w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6150w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6158w6159w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6158w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6166w6167w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6166w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6174w6175w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6174w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6182w6183w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6182w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5966w5967w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range5966w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6190w6191w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6190w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6198w6199w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6198w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5974w5975w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range5974w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5982w5983w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range5982w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5990w5991w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range5990w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5998w5999w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range5998w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6006w6007w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6006w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6014w6015w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6014w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6022w6023w(0) <= NOT wire_ccc_cordic_m_w_atannode_7_w_range6022w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6715w6716w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6715w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6796w6797w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6796w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6804w6805w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6804w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6812w6813w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6812w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6820w6821w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6820w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6828w6829w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6828w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6836w6837w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6836w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6844w6845w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6844w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6852w6853w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6852w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6860w6861w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6860w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6868w6869w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6868w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6724w6725w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6724w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6876w6877w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6876w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6884w6885w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6884w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6892w6893w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6892w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6900w6901w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6900w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6908w6909w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6908w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6916w6917w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6916w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6924w6925w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6924w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6932w6933w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6932w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6940w6941w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6940w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6948w6949w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6948w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6732w6733w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6732w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6956w6957w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6956w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6964w6965w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6964w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6740w6741w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6740w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6748w6749w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6748w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6756w6757w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6756w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6764w6765w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6764w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6772w6773w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6772w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6780w6781w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6780w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6788w6789w(0) <= NOT wire_ccc_cordic_m_w_atannode_8_w_range6788w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7476w7477w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7476w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7557w7558w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7557w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7565w7566w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7565w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7573w7574w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7573w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7581w7582w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7581w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7589w7590w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7589w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7597w7598w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7597w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7605w7606w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7605w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7613w7614w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7613w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7621w7622w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7621w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7629w7630w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7629w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7485w7486w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7485w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7637w7638w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7637w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7645w7646w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7645w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7653w7654w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7653w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7661w7662w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7661w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7669w7670w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7669w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7677w7678w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7677w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7685w7686w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7685w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7693w7694w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7693w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7701w7702w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7701w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7709w7710w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7709w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7493w7494w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7493w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7717w7718w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7717w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7725w7726w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7725w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7501w7502w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7501w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7509w7510w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7509w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7517w7518w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7517w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7525w7526w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7525w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7533w7534w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7533w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7541w7542w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7541w(0);
	wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7549w7550w(0) <= NOT wire_ccc_cordic_m_w_atannode_9_w_range7549w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range9996w9997w9998w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range9996w9997w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range9993w9994w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10033w10050w10051w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10033w10050w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10048w10049w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10038w10055w10056w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10038w10055w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10053w10054w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10043w10060w10061w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10043w10060w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10058w10059w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10048w10065w10066w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10048w10065w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10063w10064w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10053w10070w10071w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10053w10070w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10068w10069w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10058w10075w10076w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10058w10075w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10073w10074w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10063w10080w10081w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10063w10080w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10078w10079w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10068w10085w10086w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10068w10085w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10083w10084w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10073w10090w10091w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10073w10090w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10088w10089w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10078w10095w10096w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10078w10095w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10093w10094w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10003w10004w10005w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10003w10004w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10001w10002w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10083w10100w10101w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10083w10100w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10098w10099w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10088w10105w10106w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10088w10105w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10103w10104w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10093w10110w10111w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10093w10110w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10108w10109w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10098w10115w10116w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10098w10115w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10113w10114w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10103w10120w10121w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10103w10120w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10118w10119w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10108w10125w10126w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10108w10125w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10123w10124w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10113w10130w10131w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10113w10130w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10128w10129w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10118w10135w10136w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10118w10135w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10133w10134w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10123w10140w10141w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10123w10140w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10138w10139w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10128w10143w10144w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10128w10143w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10138w10139w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10009w10010w10011w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10009w10010w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10007w10008w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10133w10146w10147w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10133w10146w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10138w10139w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10138w10149w10150w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10138w10149w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10138w10139w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range9993w10015w10016w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range9993w10015w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10013w10014w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10001w10020w10021w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10001w10020w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10018w10019w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10007w10025w10026w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10007w10025w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10023w10024w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10013w10030w10031w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10013w10030w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10028w10029w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10018w10035w10036w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10018w10035w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10033w10034w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10023w10040w10041w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10023w10040w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10038w10039w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10028w10045w10046w(0) <= wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10028w10045w(0) OR wire_ccc_cordic_m_w_lg_w_pre_estimate_w_range10043w10044w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range335w338w339w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range335w338w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range320w337w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range340w343w344w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range340w343w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range325w342w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range345w348w349w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range345w348w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range330w347w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range350w353w354w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range350w353w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range335w352w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range355w358w359w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range355w358w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range340w357w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range360w363w364w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range360w363w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range345w362w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range365w368w369w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range365w368w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range350w367w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range370w373w374w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range370w373w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range355w372w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range375w378w379w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range375w378w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range360w377w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range380w383w384w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range380w383w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range365w382w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range385w388w389w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range385w388w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range370w387w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range390w393w394w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range390w393w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range375w392w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range395w398w399w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range395w398w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range380w397w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range400w403w404w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range400w403w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range385w402w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range405w408w409w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range405w408w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range390w407w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range410w413w414w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range410w413w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range395w412w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range415w418w419w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range415w418w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range400w417w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range420w423w424w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range420w423w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range405w422w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range425w428w429w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range425w428w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range410w427w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range430w433w434w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range430w433w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range415w432w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range435w438w439w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range435w438w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range420w437w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range440w443w444w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range440w443w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range425w442w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range300w303w304w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range300w303w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range289w302w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range305w308w309w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range305w308w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range294w307w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range310w313w314w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range310w313w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range297w312w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range315w318w319w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range315w318w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range300w317w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range320w323w324w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range320w323w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range305w322w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range325w328w329w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range325w328w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range310w327w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_radians_range330w333w334w(0) <= wire_ccc_cordic_m_w_lg_w_radians_range330w333w(0) OR wire_ccc_cordic_m_w_lg_w_radians_range315w332w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7019w7212w7213w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7019w7212w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7151w7210w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7078w7294w7295w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7078w7294w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7180w7293w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7084w7302w7303w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7084w7302w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7183w7301w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7090w7310w7311w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7090w7310w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7186w7309w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7096w7318w7319w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7096w7318w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7189w7317w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7102w7326w7327w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7102w7326w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7192w7325w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7108w7334w7335w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7108w7334w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7195w7333w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7114w7342w7343w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7114w7342w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7198w7341w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7120w7350w7351w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7120w7350w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7201w7349w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7126w7358w7359w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7126w7358w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7204w7357w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7132w7366w7367w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7132w7366w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7207w7365w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7024w7222w7223w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7024w7222w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7153w7221w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7138w7374w7375w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7138w7374w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range6991w7373w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7144w7382w7383w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7144w7382w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range6995w7381w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7148w7390w7391w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7148w7390w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range6997w7389w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6970w7398w7399w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6970w7398w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range6999w7397w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6975w7406w7407w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6975w7406w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7001w7405w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6977w7414w7415w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6977w7414w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7003w7413w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6979w7422w7423w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6979w7422w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7005w7421w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6981w7430w7431w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6981w7430w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7007w7429w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6983w7438w7439w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6983w7438w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7009w7437w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6985w7446w7447w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6985w7446w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7011w7445w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7030w7230w7231w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7030w7230w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7156w7229w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6987w7454w7455w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6987w7454w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7013w7453w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6989w7462w7463w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range6989w7462w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7015w7461w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7036w7238w7239w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7036w7238w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7159w7237w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7042w7246w7247w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7042w7246w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7162w7245w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7048w7254w7255w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7048w7254w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7165w7253w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7054w7262w7263w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7054w7262w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7168w7261w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7060w7270w7271w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7060w7270w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7171w7269w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7066w7278w7279w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7066w7278w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7174w7277w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7072w7286w7287w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_10_w_range7072w7286w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_10_w_range7177w7285w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7784w7968w7969w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7784w7968w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7910w7966w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7843w8050w8051w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7843w8050w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7939w8049w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7849w8058w8059w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7849w8058w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7942w8057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7855w8066w8067w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7855w8066w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7945w8065w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7861w8074w8075w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7861w8074w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7948w8073w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7867w8082w8083w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7867w8082w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7951w8081w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7873w8090w8091w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7873w8090w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7954w8089w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7879w8098w8099w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7879w8098w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7957w8097w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7885w8106w8107w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7885w8106w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7960w8105w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7891w8114w8115w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7891w8114w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7963w8113w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7897w8122w8123w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7897w8122w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7754w8121w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7789w7978w7979w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7789w7978w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7912w7977w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7903w8130w8131w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7903w8130w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7758w8129w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7907w8138w8139w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7907w8138w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7760w8137w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7731w8146w8147w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7731w8146w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7762w8145w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7736w8154w8155w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7736w8154w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7764w8153w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7738w8162w8163w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7738w8162w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7766w8161w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7740w8170w8171w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7740w8170w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7768w8169w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7742w8178w8179w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7742w8178w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7770w8177w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7744w8186w8187w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7744w8186w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7772w8185w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7746w8194w8195w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7746w8194w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7774w8193w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7748w8202w8203w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7748w8202w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7776w8201w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7795w7986w7987w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7795w7986w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7915w7985w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7750w8210w8211w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7750w8210w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7778w8209w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7752w8218w8219w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7752w8218w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7780w8217w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7801w7994w7995w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7801w7994w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7918w7993w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7807w8002w8003w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7807w8002w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7921w8001w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7813w8010w8011w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7813w8010w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7924w8009w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7819w8018w8019w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7819w8018w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7927w8017w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7825w8026w8027w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7825w8026w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7930w8025w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7831w8034w8035w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7831w8034w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7933w8033w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7837w8042w8043w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_11_w_range7837w8042w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_11_w_range7936w8041w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8544w8719w8720w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8544w8719w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8664w8717w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8603w8801w8802w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8603w8801w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8693w8800w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8609w8809w8810w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8609w8809w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8696w8808w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8615w8817w8818w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8615w8817w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8699w8816w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8621w8825w8826w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8621w8825w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8702w8824w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8627w8833w8834w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8627w8833w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8705w8832w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8633w8841w8842w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8633w8841w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8708w8840w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8639w8849w8850w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8639w8849w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8711w8848w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8645w8857w8858w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8645w8857w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8714w8856w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8651w8865w8866w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8651w8865w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8512w8864w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8657w8873w8874w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8657w8873w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8516w8872w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8549w8729w8730w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8549w8729w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8666w8728w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8661w8881w8882w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8661w8881w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8518w8880w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8487w8889w8890w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8487w8889w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8520w8888w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8492w8897w8898w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8492w8897w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8522w8896w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8494w8905w8906w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8494w8905w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8524w8904w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8496w8913w8914w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8496w8913w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8526w8912w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8498w8921w8922w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8498w8921w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8528w8920w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8500w8929w8930w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8500w8929w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8530w8928w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8502w8937w8938w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8502w8937w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8532w8936w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8504w8945w8946w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8504w8945w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8534w8944w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8506w8953w8954w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8506w8953w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8536w8952w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8555w8737w8738w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8555w8737w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8669w8736w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8508w8961w8962w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8508w8961w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8538w8960w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8510w8969w8970w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8510w8969w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8540w8968w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8561w8745w8746w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8561w8745w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8672w8744w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8567w8753w8754w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8567w8753w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8675w8752w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8573w8761w8762w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8573w8761w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8678w8760w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8579w8769w8770w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8579w8769w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8681w8768w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8585w8777w8778w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8585w8777w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8684w8776w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8591w8785w8786w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8591w8785w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8687w8784w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8597w8793w8794w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_12_w_range8597w8793w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_12_w_range8690w8792w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9299w9465w9466w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9299w9465w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9413w9463w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9358w9547w9548w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9358w9547w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9442w9546w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9364w9555w9556w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9364w9555w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9445w9554w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9370w9563w9564w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9370w9563w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9448w9562w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9376w9571w9572w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9376w9571w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9451w9570w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9382w9579w9580w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9382w9579w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9454w9578w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9388w9587w9588w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9388w9587w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9457w9586w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9394w9595w9596w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9394w9595w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9460w9594w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9400w9603w9604w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9400w9603w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9265w9602w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9406w9611w9612w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9406w9611w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9269w9610w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9410w9619w9620w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9410w9619w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9271w9618w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9304w9475w9476w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9304w9475w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9415w9474w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9238w9627w9628w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9238w9627w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9273w9626w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9243w9635w9636w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9243w9635w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9275w9634w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9245w9643w9644w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9245w9643w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9277w9642w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9247w9651w9652w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9247w9651w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9279w9650w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9249w9659w9660w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9249w9659w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9281w9658w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9251w9667w9668w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9251w9667w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9283w9666w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9253w9675w9676w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9253w9675w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9285w9674w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9255w9683w9684w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9255w9683w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9287w9682w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9257w9691w9692w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9257w9691w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9289w9690w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9259w9699w9700w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9259w9699w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9291w9698w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9310w9483w9484w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9310w9483w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9418w9482w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9261w9707w9708w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9261w9707w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9293w9706w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9263w9715w9716w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9263w9715w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9295w9714w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9316w9491w9492w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9316w9491w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9421w9490w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9322w9499w9500w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9322w9499w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9424w9498w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9328w9507w9508w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9328w9507w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9427w9506w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9334w9515w9516w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9334w9515w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9430w9514w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9340w9523w9524w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9340w9523w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9433w9522w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9346w9531w9532w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9346w9531w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9436w9530w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9352w9539w9540w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_13_w_range9352w9539w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_13_w_range9439w9538w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range719w984w985w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range719w984w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range899w982w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range778w1066w1067w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range778w1066w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range928w1065w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range784w1074w1075w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range784w1074w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range931w1073w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range790w1082w1083w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range790w1082w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range934w1081w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range796w1090w1091w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range796w1090w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range937w1089w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range802w1098w1099w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range802w1098w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range940w1097w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range808w1106w1107w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range808w1106w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range943w1105w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range814w1114w1115w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range814w1114w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range946w1113w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range820w1122w1123w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range820w1122w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range949w1121w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range826w1130w1131w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range826w1130w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range952w1129w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range832w1138w1139w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range832w1138w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range955w1137w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range724w994w995w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range724w994w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range901w993w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range838w1146w1147w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range838w1146w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range958w1145w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range844w1154w1155w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range844w1154w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range961w1153w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range850w1162w1163w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range850w1162w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range964w1161w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range856w1170w1171w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range856w1170w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range967w1169w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range862w1178w1179w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range862w1178w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range970w1177w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range868w1186w1187w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range868w1186w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range973w1185w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range874w1194w1195w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range874w1194w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range976w1193w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range880w1202w1203w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range880w1202w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range979w1201w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range886w1210w1211w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range886w1210w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range707w1209w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range892w1218w1219w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range892w1218w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range711w1217w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range730w1002w1003w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range730w1002w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range904w1001w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range896w1226w1227w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range896w1226w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range713w1225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range702w1234w1235w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range702w1234w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range715w1233w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range736w1010w1011w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range736w1010w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range907w1009w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range742w1018w1019w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range742w1018w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range910w1017w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range748w1026w1027w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range748w1026w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range913w1025w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range754w1034w1035w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range754w1034w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range916w1033w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range760w1042w1043w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range760w1042w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range919w1041w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range766w1050w1051w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range766w1050w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range922w1049w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range772w1058w1059w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_2_w_range772w1058w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_2_w_range925w1057w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1524w1780w1781w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1524w1780w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1698w1778w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1583w1862w1863w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1583w1862w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1727w1861w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1589w1870w1871w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1589w1870w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1730w1869w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1595w1878w1879w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1595w1878w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1733w1877w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1601w1886w1887w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1601w1886w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1736w1885w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1607w1894w1895w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1607w1894w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1739w1893w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1613w1902w1903w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1613w1902w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1742w1901w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1619w1910w1911w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1619w1910w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1745w1909w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1625w1918w1919w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1625w1918w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1748w1917w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1631w1926w1927w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1631w1926w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1751w1925w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1637w1934w1935w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1637w1934w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1754w1933w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1529w1790w1791w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1529w1790w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1700w1789w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1643w1942w1943w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1643w1942w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1757w1941w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1649w1950w1951w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1649w1950w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1760w1949w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1655w1958w1959w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1655w1958w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1763w1957w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1661w1966w1967w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1661w1966w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1766w1965w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1667w1974w1975w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1667w1974w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1769w1973w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1673w1982w1983w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1673w1982w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1772w1981w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1679w1990w1991w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1679w1990w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1775w1989w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1685w1998w1999w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1685w1998w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1510w1997w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1691w2006w2007w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1691w2006w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1514w2005w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1695w2014w2015w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1695w2014w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1516w2013w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1535w1798w1799w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1535w1798w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1703w1797w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1503w2022w2023w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1503w2022w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1518w2021w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1508w2030w2031w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1508w2030w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1520w2029w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1541w1806w1807w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1541w1806w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1706w1805w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1547w1814w1815w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1547w1814w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1709w1813w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1553w1822w1823w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1553w1822w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1712w1821w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1559w1830w1831w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1559w1830w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1715w1829w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1565w1838w1839w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1565w1838w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1718w1837w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1571w1846w1847w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1571w1846w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1721w1845w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1577w1854w1855w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_3_w_range1577w1854w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_3_w_range1724w1853w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2324w2571w2572w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2324w2571w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2492w2569w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2383w2653w2654w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2383w2653w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2521w2652w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2389w2661w2662w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2389w2661w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2524w2660w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2395w2669w2670w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2395w2669w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2527w2668w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2401w2677w2678w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2401w2677w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2530w2676w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2407w2685w2686w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2407w2685w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2533w2684w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2413w2693w2694w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2413w2693w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2536w2692w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2419w2701w2702w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2419w2701w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2539w2700w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2425w2709w2710w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2425w2709w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2542w2708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2431w2717w2718w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2431w2717w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2545w2716w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2437w2725w2726w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2437w2725w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2548w2724w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2329w2581w2582w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2329w2581w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2494w2580w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2443w2733w2734w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2443w2733w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2551w2732w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2449w2741w2742w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2449w2741w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2554w2740w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2455w2749w2750w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2455w2749w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2557w2748w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2461w2757w2758w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2461w2757w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2560w2756w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2467w2765w2766w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2467w2765w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2563w2764w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2473w2773w2774w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2473w2773w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2566w2772w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2479w2781w2782w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2479w2781w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2308w2780w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2485w2789w2790w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2485w2789w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2312w2788w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2489w2797w2798w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2489w2797w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2314w2796w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2299w2805w2806w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2299w2805w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2316w2804w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2335w2589w2590w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2335w2589w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2497w2588w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2304w2813w2814w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2304w2813w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2318w2812w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2306w2821w2822w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2306w2821w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2320w2820w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2341w2597w2598w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2341w2597w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2500w2596w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2347w2605w2606w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2347w2605w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2503w2604w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2353w2613w2614w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2353w2613w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2506w2612w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2359w2621w2622w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2359w2621w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2509w2620w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2365w2629w2630w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2365w2629w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2512w2628w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2371w2637w2638w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2371w2637w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2515w2636w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2377w2645w2646w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_4_w_range2377w2645w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_4_w_range2518w2644w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3119w3357w3358w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3119w3357w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3281w3355w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3178w3439w3440w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3178w3439w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3310w3438w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3184w3447w3448w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3184w3447w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3313w3446w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3190w3455w3456w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3190w3455w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3316w3454w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3196w3463w3464w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3196w3463w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3319w3462w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3202w3471w3472w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3202w3471w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3322w3470w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3208w3479w3480w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3208w3479w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3325w3478w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3214w3487w3488w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3214w3487w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3328w3486w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3220w3495w3496w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3220w3495w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3331w3494w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3226w3503w3504w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3226w3503w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3334w3502w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3232w3511w3512w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3232w3511w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3337w3510w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3124w3367w3368w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3124w3367w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3283w3366w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3238w3519w3520w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3238w3519w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3340w3518w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3244w3527w3528w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3244w3527w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3343w3526w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3250w3535w3536w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3250w3535w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3346w3534w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3256w3543w3544w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3256w3543w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3349w3542w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3262w3551w3552w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3262w3551w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3352w3550w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3268w3559w3560w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3268w3559w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3101w3558w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3274w3567w3568w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3274w3567w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3105w3566w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3278w3575w3576w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3278w3575w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3107w3574w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3090w3583w3584w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3090w3583w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3109w3582w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3095w3591w3592w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3095w3591w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3111w3590w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3130w3375w3376w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3130w3375w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3286w3374w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3097w3599w3600w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3097w3599w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3113w3598w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3099w3607w3608w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3099w3607w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3115w3606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3136w3383w3384w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3136w3383w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3289w3382w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3142w3391w3392w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3142w3391w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3292w3390w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3148w3399w3400w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3148w3399w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3295w3398w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3154w3407w3408w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3154w3407w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3298w3406w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3160w3415w3416w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3160w3415w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3301w3414w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3166w3423w3424w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3166w3423w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3304w3422w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3172w3431w3432w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_5_w_range3172w3431w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_5_w_range3307w3430w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3909w4138w4139w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3909w4138w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4065w4136w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3968w4220w4221w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3968w4220w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4094w4219w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3974w4228w4229w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3974w4228w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4097w4227w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3980w4236w4237w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3980w4236w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4100w4235w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3986w4244w4245w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3986w4244w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4103w4243w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3992w4252w4253w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3992w4252w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4106w4251w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3998w4260w4261w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3998w4260w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4109w4259w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4004w4268w4269w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4004w4268w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4112w4267w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4010w4276w4277w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4010w4276w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4115w4275w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4016w4284w4285w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4016w4284w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4118w4283w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4022w4292w4293w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4022w4292w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4121w4291w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3914w4148w4149w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3914w4148w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4067w4147w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4028w4300w4301w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4028w4300w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4124w4299w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4034w4308w4309w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4034w4308w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4127w4307w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4040w4316w4317w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4040w4316w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4130w4315w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4046w4324w4325w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4046w4324w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4133w4323w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4052w4332w4333w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4052w4332w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3889w4331w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4058w4340w4341w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4058w4340w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3893w4339w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4062w4348w4349w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range4062w4348w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3895w4347w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3876w4356w4357w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3876w4356w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3897w4355w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3881w4364w4365w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3881w4364w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3899w4363w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3883w4372w4373w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3883w4372w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3901w4371w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3920w4156w4157w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3920w4156w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4070w4155w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3885w4380w4381w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3885w4380w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3903w4379w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3887w4388w4389w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3887w4388w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range3905w4387w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3926w4164w4165w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3926w4164w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4073w4163w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3932w4172w4173w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3932w4172w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4076w4171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3938w4180w4181w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3938w4180w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4079w4179w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3944w4188w4189w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3944w4188w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4082w4187w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3950w4196w4197w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3950w4196w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4085w4195w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3956w4204w4205w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3956w4204w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4088w4203w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3962w4212w4213w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_6_w_range3962w4212w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_6_w_range4091w4211w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4694w4914w4915w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4694w4914w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4844w4912w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4753w4996w4997w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4753w4996w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4873w4995w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4759w5004w5005w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4759w5004w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4876w5003w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4765w5012w5013w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4765w5012w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4879w5011w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4771w5020w5021w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4771w5020w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4882w5019w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4777w5028w5029w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4777w5028w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4885w5027w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4783w5036w5037w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4783w5036w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4888w5035w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4789w5044w5045w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4789w5044w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4891w5043w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4795w5052w5053w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4795w5052w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4894w5051w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4801w5060w5061w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4801w5060w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4897w5059w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4807w5068w5069w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4807w5068w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4900w5067w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4699w4924w4925w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4699w4924w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4846w4923w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4813w5076w5077w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4813w5076w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4903w5075w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4819w5084w5085w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4819w5084w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4906w5083w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4825w5092w5093w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4825w5092w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4909w5091w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4831w5100w5101w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4831w5100w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4672w5099w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4837w5108w5109w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4837w5108w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4676w5107w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4841w5116w5117w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4841w5116w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4678w5115w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4657w5124w5125w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4657w5124w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4680w5123w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4662w5132w5133w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4662w5132w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4682w5131w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4664w5140w5141w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4664w5140w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4684w5139w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4666w5148w5149w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4666w5148w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4686w5147w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4705w4932w4933w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4705w4932w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4849w4931w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4668w5156w5157w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4668w5156w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4688w5155w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4670w5164w5165w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4670w5164w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4690w5163w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4711w4940w4941w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4711w4940w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4852w4939w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4717w4948w4949w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4717w4948w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4855w4947w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4723w4956w4957w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4723w4956w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4858w4955w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4729w4964w4965w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4729w4964w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4861w4963w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4735w4972w4973w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4735w4972w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4864w4971w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4741w4980w4981w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4741w4980w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4867w4979w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4747w4988w4989w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_7_w_range4747w4988w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_7_w_range4870w4987w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5474w5685w5686w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5474w5685w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5618w5683w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5533w5767w5768w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5533w5767w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5647w5766w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5539w5775w5776w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5539w5775w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5650w5774w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5545w5783w5784w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5545w5783w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5653w5782w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5551w5791w5792w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5551w5791w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5656w5790w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5557w5799w5800w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5557w5799w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5659w5798w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5563w5807w5808w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5563w5807w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5662w5806w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5569w5815w5816w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5569w5815w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5665w5814w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5575w5823w5824w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5575w5823w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5668w5822w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5581w5831w5832w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5581w5831w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5671w5830w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5587w5839w5840w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5587w5839w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5674w5838w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5479w5695w5696w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5479w5695w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5620w5694w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5593w5847w5848w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5593w5847w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5677w5846w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5599w5855w5856w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5599w5855w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5680w5854w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5605w5863w5864w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5605w5863w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5450w5862w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5611w5871w5872w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5611w5871w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5454w5870w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5615w5879w5880w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5615w5879w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5456w5878w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5433w5887w5888w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5433w5887w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5458w5886w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5438w5895w5896w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5438w5895w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5460w5894w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5440w5903w5904w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5440w5903w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5462w5902w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5442w5911w5912w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5442w5911w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5464w5910w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5444w5919w5920w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5444w5919w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5466w5918w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5485w5703w5704w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5485w5703w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5623w5702w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5446w5927w5928w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5446w5927w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5468w5926w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5448w5935w5936w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5448w5935w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5470w5934w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5491w5711w5712w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5491w5711w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5626w5710w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5497w5719w5720w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5497w5719w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5629w5718w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5503w5727w5728w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5503w5727w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5632w5726w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5509w5735w5736w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5509w5735w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5635w5734w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5515w5743w5744w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5515w5743w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5638w5742w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5521w5751w5752w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5521w5751w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5641w5750w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5527w5759w5760w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_8_w_range5527w5759w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_8_w_range5644w5758w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6249w6451w6452w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6249w6451w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6387w6449w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6308w6533w6534w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6308w6533w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6416w6532w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6314w6541w6542w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6314w6541w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6419w6540w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6320w6549w6550w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6320w6549w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6422w6548w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6326w6557w6558w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6326w6557w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6425w6556w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6332w6565w6566w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6332w6565w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6428w6564w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6338w6573w6574w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6338w6573w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6431w6572w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6344w6581w6582w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6344w6581w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6434w6580w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6350w6589w6590w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6350w6589w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6437w6588w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6356w6597w6598w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6356w6597w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6440w6596w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6362w6605w6606w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6362w6605w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6443w6604w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6254w6461w6462w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6254w6461w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6389w6460w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6368w6613w6614w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6368w6613w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6446w6612w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6374w6621w6622w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6374w6621w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6223w6620w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6380w6629w6630w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6380w6629w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6227w6628w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6384w6637w6638w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6384w6637w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6229w6636w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6204w6645w6646w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6204w6645w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6231w6644w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6209w6653w6654w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6209w6653w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6233w6652w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6211w6661w6662w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6211w6661w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6235w6660w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6213w6669w6670w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6213w6669w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6237w6668w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6215w6677w6678w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6215w6677w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6239w6676w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6217w6685w6686w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6217w6685w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6241w6684w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6260w6469w6470w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6260w6469w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6392w6468w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6219w6693w6694w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6219w6693w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6243w6692w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6221w6701w6702w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6221w6701w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6245w6700w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6266w6477w6478w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6266w6477w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6395w6476w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6272w6485w6486w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6272w6485w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6398w6484w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6278w6493w6494w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6278w6493w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6401w6492w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6284w6501w6502w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6284w6501w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6404w6500w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6290w6509w6510w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6290w6509w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6407w6508w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6296w6517w6518w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6296w6517w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6410w6516w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6302w6525w6526w(0) <= wire_ccc_cordic_m_w_lg_w_x_prenodeone_9_w_range6302w6525w(0) OR wire_ccc_cordic_m_w_lg_w_x_prenodetwo_9_w_range6413w6524w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7021w7217w7218w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7021w7217w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7152w7216w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7080w7298w7299w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7080w7298w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7181w7297w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7086w7306w7307w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7086w7306w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7184w7305w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7092w7314w7315w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7092w7314w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7187w7313w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7098w7322w7323w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7098w7322w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7190w7321w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7104w7330w7331w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7104w7330w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7193w7329w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7110w7338w7339w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7110w7338w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7196w7337w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7116w7346w7347w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7116w7346w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7199w7345w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7122w7354w7355w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7122w7354w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7202w7353w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7128w7362w7363w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7128w7362w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7205w7361w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7134w7370w7371w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7134w7370w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7208w7369w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7026w7226w7227w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7026w7226w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7154w7225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7140w7378w7379w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7140w7378w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range6993w7377w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7146w7386w7387w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7146w7386w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range6996w7385w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7149w7394w7395w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7149w7394w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range6998w7393w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6973w7402w7403w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6973w7402w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7000w7401w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6976w7410w7411w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6976w7410w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7002w7409w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6978w7418w7419w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6978w7418w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7004w7417w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6980w7426w7427w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6980w7426w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7006w7425w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6982w7434w7435w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6982w7434w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7008w7433w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6984w7442w7443w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6984w7442w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7010w7441w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6986w7450w7451w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6986w7450w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7012w7449w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7032w7234w7235w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7032w7234w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7157w7233w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6988w7458w7459w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6988w7458w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7014w7457w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6990w7466w7467w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range6990w7466w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7016w7465w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7038w7242w7243w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7038w7242w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7160w7241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7044w7250w7251w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7044w7250w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7163w7249w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7050w7258w7259w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7050w7258w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7166w7257w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7056w7266w7267w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7056w7266w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7169w7265w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7062w7274w7275w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7062w7274w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7172w7273w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7068w7282w7283w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7068w7282w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7175w7281w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7074w7290w7291w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_10_w_range7074w7290w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_10_w_range7178w7289w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7786w7973w7974w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7786w7973w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7911w7972w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7845w8054w8055w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7845w8054w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7940w8053w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7851w8062w8063w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7851w8062w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7943w8061w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7857w8070w8071w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7857w8070w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7946w8069w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7863w8078w8079w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7863w8078w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7949w8077w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7869w8086w8087w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7869w8086w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7952w8085w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7875w8094w8095w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7875w8094w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7955w8093w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7881w8102w8103w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7881w8102w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7958w8101w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7887w8110w8111w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7887w8110w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7961w8109w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7893w8118w8119w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7893w8118w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7964w8117w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7899w8126w8127w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7899w8126w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7756w8125w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7791w7982w7983w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7791w7982w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7913w7981w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7905w8134w8135w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7905w8134w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7759w8133w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7908w8142w8143w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7908w8142w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7761w8141w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7734w8150w8151w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7734w8150w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7763w8149w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7737w8158w8159w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7737w8158w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7765w8157w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7739w8166w8167w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7739w8166w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7767w8165w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7741w8174w8175w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7741w8174w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7769w8173w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7743w8182w8183w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7743w8182w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7771w8181w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7745w8190w8191w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7745w8190w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7773w8189w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7747w8198w8199w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7747w8198w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7775w8197w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7749w8206w8207w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7749w8206w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7777w8205w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7797w7990w7991w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7797w7990w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7916w7989w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7751w8214w8215w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7751w8214w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7779w8213w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7753w8222w8223w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7753w8222w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7781w8221w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7803w7998w7999w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7803w7998w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7919w7997w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7809w8006w8007w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7809w8006w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7922w8005w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7815w8014w8015w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7815w8014w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7925w8013w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7821w8022w8023w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7821w8022w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7928w8021w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7827w8030w8031w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7827w8030w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7931w8029w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7833w8038w8039w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7833w8038w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7934w8037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7839w8046w8047w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_11_w_range7839w8046w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_11_w_range7937w8045w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8546w8724w8725w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8546w8724w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8665w8723w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8605w8805w8806w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8605w8805w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8694w8804w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8611w8813w8814w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8611w8813w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8697w8812w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8617w8821w8822w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8617w8821w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8700w8820w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8623w8829w8830w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8623w8829w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8703w8828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8629w8837w8838w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8629w8837w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8706w8836w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8635w8845w8846w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8635w8845w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8709w8844w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8641w8853w8854w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8641w8853w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8712w8852w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8647w8861w8862w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8647w8861w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8715w8860w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8653w8869w8870w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8653w8869w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8514w8868w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8659w8877w8878w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8659w8877w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8517w8876w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8551w8733w8734w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8551w8733w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8667w8732w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8662w8885w8886w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8662w8885w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8519w8884w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8490w8893w8894w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8490w8893w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8521w8892w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8493w8901w8902w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8493w8901w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8523w8900w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8495w8909w8910w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8495w8909w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8525w8908w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8497w8917w8918w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8497w8917w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8527w8916w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8499w8925w8926w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8499w8925w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8529w8924w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8501w8933w8934w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8501w8933w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8531w8932w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8503w8941w8942w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8503w8941w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8533w8940w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8505w8949w8950w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8505w8949w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8535w8948w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8507w8957w8958w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8507w8957w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8537w8956w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8557w8741w8742w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8557w8741w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8670w8740w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8509w8965w8966w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8509w8965w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8539w8964w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8511w8973w8974w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8511w8973w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8541w8972w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8563w8749w8750w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8563w8749w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8673w8748w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8569w8757w8758w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8569w8757w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8676w8756w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8575w8765w8766w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8575w8765w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8679w8764w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8581w8773w8774w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8581w8773w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8682w8772w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8587w8781w8782w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8587w8781w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8685w8780w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8593w8789w8790w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8593w8789w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8688w8788w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8599w8797w8798w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_12_w_range8599w8797w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_12_w_range8691w8796w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9301w9470w9471w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9301w9470w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9414w9469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9360w9551w9552w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9360w9551w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9443w9550w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9366w9559w9560w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9366w9559w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9446w9558w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9372w9567w9568w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9372w9567w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9449w9566w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9378w9575w9576w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9378w9575w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9452w9574w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9384w9583w9584w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9384w9583w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9455w9582w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9390w9591w9592w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9390w9591w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9458w9590w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9396w9599w9600w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9396w9599w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9461w9598w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9402w9607w9608w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9402w9607w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9267w9606w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9408w9615w9616w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9408w9615w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9270w9614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9411w9623w9624w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9411w9623w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9272w9622w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9306w9479w9480w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9306w9479w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9416w9478w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9241w9631w9632w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9241w9631w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9274w9630w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9244w9639w9640w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9244w9639w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9276w9638w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9246w9647w9648w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9246w9647w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9278w9646w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9248w9655w9656w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9248w9655w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9280w9654w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9250w9663w9664w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9250w9663w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9282w9662w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9252w9671w9672w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9252w9671w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9284w9670w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9254w9679w9680w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9254w9679w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9286w9678w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9256w9687w9688w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9256w9687w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9288w9686w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9258w9695w9696w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9258w9695w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9290w9694w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9260w9703w9704w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9260w9703w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9292w9702w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9312w9487w9488w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9312w9487w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9419w9486w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9262w9711w9712w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9262w9711w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9294w9710w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9264w9719w9720w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9264w9719w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9296w9718w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9318w9495w9496w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9318w9495w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9422w9494w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9324w9503w9504w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9324w9503w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9425w9502w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9330w9511w9512w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9330w9511w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9428w9510w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9336w9519w9520w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9336w9519w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9431w9518w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9342w9527w9528w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9342w9527w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9434w9526w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9348w9535w9536w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9348w9535w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9437w9534w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9354w9543w9544w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_13_w_range9354w9543w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_13_w_range9440w9542w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range721w989w990w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range721w989w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range900w988w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range780w1070w1071w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range780w1070w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range929w1069w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range786w1078w1079w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range786w1078w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range932w1077w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range792w1086w1087w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range792w1086w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range935w1085w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range798w1094w1095w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range798w1094w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range938w1093w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range804w1102w1103w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range804w1102w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range941w1101w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range810w1110w1111w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range810w1110w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range944w1109w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range816w1118w1119w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range816w1118w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range947w1117w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range822w1126w1127w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range822w1126w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range950w1125w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range828w1134w1135w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range828w1134w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range953w1133w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range834w1142w1143w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range834w1142w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range956w1141w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range726w998w999w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range726w998w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range902w997w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range840w1150w1151w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range840w1150w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range959w1149w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range846w1158w1159w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range846w1158w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range962w1157w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range852w1166w1167w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range852w1166w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range965w1165w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range858w1174w1175w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range858w1174w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range968w1173w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range864w1182w1183w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range864w1182w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range971w1181w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range870w1190w1191w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range870w1190w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range974w1189w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range876w1198w1199w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range876w1198w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range977w1197w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range882w1206w1207w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range882w1206w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range980w1205w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range888w1214w1215w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range888w1214w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range709w1213w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range894w1222w1223w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range894w1222w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range712w1221w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range732w1006w1007w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range732w1006w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range905w1005w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range897w1230w1231w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range897w1230w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range714w1229w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range705w1238w1239w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range705w1238w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range716w1237w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range738w1014w1015w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range738w1014w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range908w1013w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range744w1022w1023w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range744w1022w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range911w1021w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range750w1030w1031w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range750w1030w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range914w1029w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range756w1038w1039w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range756w1038w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range917w1037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range762w1046w1047w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range762w1046w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range920w1045w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range768w1054w1055w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range768w1054w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range923w1053w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range774w1062w1063w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_2_w_range774w1062w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_2_w_range926w1061w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1526w1785w1786w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1526w1785w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1699w1784w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1585w1866w1867w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1585w1866w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1728w1865w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1591w1874w1875w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1591w1874w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1731w1873w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1597w1882w1883w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1597w1882w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1734w1881w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1603w1890w1891w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1603w1890w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1737w1889w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1609w1898w1899w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1609w1898w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1740w1897w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1615w1906w1907w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1615w1906w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1743w1905w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1621w1914w1915w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1621w1914w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1746w1913w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1627w1922w1923w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1627w1922w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1749w1921w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1633w1930w1931w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1633w1930w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1752w1929w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1639w1938w1939w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1639w1938w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1755w1937w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1531w1794w1795w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1531w1794w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1701w1793w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1645w1946w1947w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1645w1946w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1758w1945w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1651w1954w1955w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1651w1954w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1761w1953w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1657w1962w1963w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1657w1962w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1764w1961w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1663w1970w1971w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1663w1970w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1767w1969w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1669w1978w1979w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1669w1978w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1770w1977w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1675w1986w1987w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1675w1986w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1773w1985w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1681w1994w1995w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1681w1994w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1776w1993w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1687w2002w2003w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1687w2002w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1512w2001w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1693w2010w2011w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1693w2010w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1515w2009w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1696w2018w2019w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1696w2018w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1517w2017w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1537w1802w1803w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1537w1802w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1704w1801w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1506w2026w2027w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1506w2026w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1519w2025w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1509w2034w2035w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1509w2034w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1521w2033w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1543w1810w1811w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1543w1810w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1707w1809w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1549w1818w1819w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1549w1818w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1710w1817w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1555w1826w1827w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1555w1826w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1713w1825w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1561w1834w1835w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1561w1834w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1716w1833w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1567w1842w1843w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1567w1842w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1719w1841w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1573w1850w1851w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1573w1850w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1722w1849w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1579w1858w1859w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_3_w_range1579w1858w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_3_w_range1725w1857w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2326w2576w2577w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2326w2576w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2493w2575w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2385w2657w2658w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2385w2657w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2522w2656w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2391w2665w2666w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2391w2665w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2525w2664w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2397w2673w2674w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2397w2673w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2528w2672w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2403w2681w2682w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2403w2681w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2531w2680w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2409w2689w2690w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2409w2689w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2534w2688w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2415w2697w2698w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2415w2697w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2537w2696w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2421w2705w2706w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2421w2705w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2540w2704w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2427w2713w2714w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2427w2713w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2543w2712w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2433w2721w2722w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2433w2721w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2546w2720w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2439w2729w2730w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2439w2729w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2549w2728w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2331w2585w2586w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2331w2585w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2495w2584w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2445w2737w2738w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2445w2737w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2552w2736w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2451w2745w2746w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2451w2745w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2555w2744w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2457w2753w2754w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2457w2753w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2558w2752w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2463w2761w2762w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2463w2761w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2561w2760w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2469w2769w2770w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2469w2769w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2564w2768w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2475w2777w2778w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2475w2777w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2567w2776w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2481w2785w2786w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2481w2785w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2310w2784w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2487w2793w2794w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2487w2793w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2313w2792w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2490w2801w2802w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2490w2801w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2315w2800w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2302w2809w2810w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2302w2809w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2317w2808w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2337w2593w2594w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2337w2593w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2498w2592w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2305w2817w2818w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2305w2817w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2319w2816w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2307w2825w2826w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2307w2825w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2321w2824w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2343w2601w2602w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2343w2601w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2501w2600w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2349w2609w2610w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2349w2609w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2504w2608w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2355w2617w2618w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2355w2617w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2507w2616w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2361w2625w2626w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2361w2625w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2510w2624w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2367w2633w2634w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2367w2633w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2513w2632w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2373w2641w2642w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2373w2641w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2516w2640w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2379w2649w2650w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_4_w_range2379w2649w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_4_w_range2519w2648w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3121w3362w3363w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3121w3362w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3282w3361w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3180w3443w3444w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3180w3443w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3311w3442w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3186w3451w3452w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3186w3451w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3314w3450w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3192w3459w3460w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3192w3459w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3317w3458w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3198w3467w3468w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3198w3467w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3320w3466w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3204w3475w3476w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3204w3475w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3323w3474w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3210w3483w3484w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3210w3483w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3326w3482w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3216w3491w3492w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3216w3491w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3329w3490w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3222w3499w3500w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3222w3499w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3332w3498w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3228w3507w3508w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3228w3507w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3335w3506w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3234w3515w3516w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3234w3515w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3338w3514w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3126w3371w3372w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3126w3371w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3284w3370w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3240w3523w3524w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3240w3523w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3341w3522w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3246w3531w3532w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3246w3531w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3344w3530w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3252w3539w3540w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3252w3539w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3347w3538w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3258w3547w3548w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3258w3547w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3350w3546w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3264w3555w3556w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3264w3555w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3353w3554w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3270w3563w3564w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3270w3563w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3103w3562w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3276w3571w3572w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3276w3571w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3106w3570w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3279w3579w3580w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3279w3579w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3108w3578w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3093w3587w3588w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3093w3587w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3110w3586w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3096w3595w3596w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3096w3595w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3112w3594w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3132w3379w3380w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3132w3379w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3287w3378w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3098w3603w3604w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3098w3603w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3114w3602w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3100w3611w3612w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3100w3611w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3116w3610w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3138w3387w3388w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3138w3387w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3290w3386w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3144w3395w3396w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3144w3395w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3293w3394w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3150w3403w3404w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3150w3403w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3296w3402w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3156w3411w3412w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3156w3411w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3299w3410w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3162w3419w3420w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3162w3419w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3302w3418w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3168w3427w3428w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3168w3427w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3305w3426w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3174w3435w3436w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_5_w_range3174w3435w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_5_w_range3308w3434w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3911w4143w4144w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3911w4143w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4066w4142w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3970w4224w4225w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3970w4224w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4095w4223w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3976w4232w4233w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3976w4232w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4098w4231w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3982w4240w4241w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3982w4240w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4101w4239w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3988w4248w4249w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3988w4248w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4104w4247w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3994w4256w4257w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3994w4256w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4107w4255w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4000w4264w4265w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4000w4264w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4110w4263w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4006w4272w4273w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4006w4272w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4113w4271w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4012w4280w4281w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4012w4280w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4116w4279w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4018w4288w4289w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4018w4288w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4119w4287w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4024w4296w4297w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4024w4296w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4122w4295w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3916w4152w4153w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3916w4152w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4068w4151w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4030w4304w4305w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4030w4304w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4125w4303w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4036w4312w4313w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4036w4312w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4128w4311w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4042w4320w4321w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4042w4320w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4131w4319w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4048w4328w4329w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4048w4328w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4134w4327w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4054w4336w4337w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4054w4336w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3891w4335w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4060w4344w4345w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4060w4344w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3894w4343w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4063w4352w4353w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range4063w4352w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3896w4351w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3879w4360w4361w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3879w4360w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3898w4359w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3882w4368w4369w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3882w4368w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3900w4367w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3884w4376w4377w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3884w4376w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3902w4375w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3922w4160w4161w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3922w4160w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4071w4159w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3886w4384w4385w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3886w4384w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3904w4383w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3888w4392w4393w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3888w4392w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range3906w4391w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3928w4168w4169w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3928w4168w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4074w4167w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3934w4176w4177w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3934w4176w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4077w4175w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3940w4184w4185w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3940w4184w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4080w4183w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3946w4192w4193w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3946w4192w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4083w4191w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3952w4200w4201w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3952w4200w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4086w4199w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3958w4208w4209w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3958w4208w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4089w4207w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3964w4216w4217w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_6_w_range3964w4216w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_6_w_range4092w4215w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4696w4919w4920w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4696w4919w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4845w4918w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4755w5000w5001w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4755w5000w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4874w4999w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4761w5008w5009w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4761w5008w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4877w5007w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4767w5016w5017w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4767w5016w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4880w5015w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4773w5024w5025w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4773w5024w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4883w5023w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4779w5032w5033w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4779w5032w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4886w5031w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4785w5040w5041w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4785w5040w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4889w5039w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4791w5048w5049w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4791w5048w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4892w5047w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4797w5056w5057w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4797w5056w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4895w5055w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4803w5064w5065w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4803w5064w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4898w5063w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4809w5072w5073w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4809w5072w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4901w5071w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4701w4928w4929w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4701w4928w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4847w4927w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4815w5080w5081w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4815w5080w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4904w5079w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4821w5088w5089w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4821w5088w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4907w5087w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4827w5096w5097w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4827w5096w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4910w5095w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4833w5104w5105w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4833w5104w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4674w5103w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4839w5112w5113w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4839w5112w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4677w5111w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4842w5120w5121w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4842w5120w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4679w5119w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4660w5128w5129w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4660w5128w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4681w5127w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4663w5136w5137w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4663w5136w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4683w5135w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4665w5144w5145w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4665w5144w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4685w5143w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4667w5152w5153w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4667w5152w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4687w5151w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4707w4936w4937w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4707w4936w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4850w4935w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4669w5160w5161w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4669w5160w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4689w5159w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4671w5168w5169w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4671w5168w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4691w5167w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4713w4944w4945w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4713w4944w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4853w4943w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4719w4952w4953w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4719w4952w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4856w4951w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4725w4960w4961w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4725w4960w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4859w4959w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4731w4968w4969w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4731w4968w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4862w4967w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4737w4976w4977w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4737w4976w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4865w4975w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4743w4984w4985w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4743w4984w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4868w4983w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4749w4992w4993w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_7_w_range4749w4992w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_7_w_range4871w4991w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5476w5690w5691w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5476w5690w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5619w5689w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5535w5771w5772w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5535w5771w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5648w5770w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5541w5779w5780w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5541w5779w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5651w5778w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5547w5787w5788w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5547w5787w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5654w5786w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5553w5795w5796w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5553w5795w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5657w5794w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5559w5803w5804w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5559w5803w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5660w5802w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5565w5811w5812w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5565w5811w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5663w5810w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5571w5819w5820w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5571w5819w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5666w5818w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5577w5827w5828w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5577w5827w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5669w5826w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5583w5835w5836w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5583w5835w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5672w5834w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5589w5843w5844w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5589w5843w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5675w5842w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5481w5699w5700w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5481w5699w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5621w5698w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5595w5851w5852w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5595w5851w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5678w5850w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5601w5859w5860w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5601w5859w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5681w5858w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5607w5867w5868w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5607w5867w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5452w5866w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5613w5875w5876w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5613w5875w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5455w5874w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5616w5883w5884w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5616w5883w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5457w5882w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5436w5891w5892w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5436w5891w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5459w5890w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5439w5899w5900w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5439w5899w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5461w5898w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5441w5907w5908w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5441w5907w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5463w5906w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5443w5915w5916w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5443w5915w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5465w5914w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5445w5923w5924w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5445w5923w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5467w5922w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5487w5707w5708w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5487w5707w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5624w5706w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5447w5931w5932w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5447w5931w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5469w5930w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5449w5939w5940w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5449w5939w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5471w5938w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5493w5715w5716w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5493w5715w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5627w5714w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5499w5723w5724w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5499w5723w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5630w5722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5505w5731w5732w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5505w5731w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5633w5730w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5511w5739w5740w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5511w5739w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5636w5738w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5517w5747w5748w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5517w5747w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5639w5746w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5523w5755w5756w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5523w5755w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5642w5754w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5529w5763w5764w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_8_w_range5529w5763w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_8_w_range5645w5762w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6251w6456w6457w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6251w6456w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6388w6455w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6310w6537w6538w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6310w6537w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6417w6536w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6316w6545w6546w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6316w6545w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6420w6544w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6322w6553w6554w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6322w6553w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6423w6552w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6328w6561w6562w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6328w6561w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6426w6560w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6334w6569w6570w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6334w6569w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6429w6568w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6340w6577w6578w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6340w6577w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6432w6576w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6346w6585w6586w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6346w6585w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6435w6584w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6352w6593w6594w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6352w6593w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6438w6592w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6358w6601w6602w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6358w6601w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6441w6600w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6364w6609w6610w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6364w6609w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6444w6608w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6256w6465w6466w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6256w6465w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6390w6464w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6370w6617w6618w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6370w6617w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6447w6616w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6376w6625w6626w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6376w6625w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6225w6624w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6382w6633w6634w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6382w6633w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6228w6632w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6385w6641w6642w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6385w6641w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6230w6640w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6207w6649w6650w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6207w6649w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6232w6648w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6210w6657w6658w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6210w6657w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6234w6656w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6212w6665w6666w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6212w6665w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6236w6664w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6214w6673w6674w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6214w6673w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6238w6672w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6216w6681w6682w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6216w6681w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6240w6680w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6218w6689w6690w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6218w6689w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6242w6688w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6262w6473w6474w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6262w6473w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6393w6472w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6220w6697w6698w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6220w6697w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6244w6696w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6222w6705w6706w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6222w6705w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6246w6704w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6268w6481w6482w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6268w6481w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6396w6480w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6274w6489w6490w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6274w6489w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6399w6488w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6280w6497w6498w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6280w6497w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6402w6496w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6286w6505w6506w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6286w6505w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6405w6504w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6292w6513w6514w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6292w6513w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6408w6512w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6298w6521w6522w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6298w6521w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6411w6520w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6304w6529w6530w(0) <= wire_ccc_cordic_m_w_lg_w_y_prenodeone_9_w_range6304w6529w(0) OR wire_ccc_cordic_m_w_lg_w_y_prenodetwo_9_w_range6414w6528w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8232w8233w8234w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8232w8233w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8313w8314w8315w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8313w8314w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8321w8322w8323w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8321w8322w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8329w8330w8331w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8329w8330w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8337w8338w8339w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8337w8338w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8345w8346w8347w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8345w8346w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8353w8354w8355w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8353w8354w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8361w8362w8363w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8361w8362w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8369w8370w8371w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8369w8370w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8377w8378w8379w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8377w8378w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8385w8386w8387w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8385w8386w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8241w8242w8243w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8241w8242w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8393w8394w8395w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8393w8394w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8401w8402w8403w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8401w8402w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8409w8410w8411w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8409w8410w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8417w8418w8419w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8417w8418w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8425w8426w8427w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8425w8426w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8433w8434w8435w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8433w8434w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8441w8442w8443w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8441w8442w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8449w8450w8451w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8449w8450w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8457w8458w8459w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8457w8458w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8465w8466w8467w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8465w8466w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8249w8250w8251w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8249w8250w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8473w8474w8475w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8473w8474w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8481w8482w8483w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8481w8482w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8257w8258w8259w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8257w8258w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8265w8266w8267w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8265w8266w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8273w8274w8275w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8273w8274w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8281w8282w8283w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8281w8282w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8289w8290w8291w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8289w8290w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8297w8298w8299w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8297w8298w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8305w8306w8307w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_10_w_range8305w8306w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range8983w8984w8985w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range8983w8984w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9064w9065w9066w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9064w9065w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9072w9073w9074w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9072w9073w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9080w9081w9082w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9080w9081w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9088w9089w9090w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9088w9089w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9096w9097w9098w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9096w9097w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9104w9105w9106w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9104w9105w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9112w9113w9114w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9112w9113w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9120w9121w9122w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9120w9121w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9128w9129w9130w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9128w9129w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9136w9137w9138w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9136w9137w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range8992w8993w8994w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range8992w8993w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9144w9145w9146w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9144w9145w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9152w9153w9154w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9152w9153w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9160w9161w9162w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9160w9161w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9168w9169w9170w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9168w9169w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9176w9177w9178w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9176w9177w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9184w9185w9186w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9184w9185w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9192w9193w9194w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9192w9193w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9200w9201w9202w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9200w9201w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9208w9209w9210w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9208w9209w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9216w9217w9218w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9216w9217w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9000w9001w9002w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9000w9001w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9224w9225w9226w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9224w9225w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9232w9233w9234w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9232w9233w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9008w9009w9010w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9008w9009w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9016w9017w9018w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9016w9017w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9024w9025w9026w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9024w9025w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9032w9033w9034w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9032w9033w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9040w9041w9042w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9040w9041w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9048w9049w9050w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9048w9049w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9056w9057w9058w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_11_w_range9056w9057w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9729w9730w9731w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9729w9730w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9810w9811w9812w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9810w9811w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9818w9819w9820w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9818w9819w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9826w9827w9828w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9826w9827w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9834w9835w9836w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9834w9835w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9842w9843w9844w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9842w9843w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9850w9851w9852w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9850w9851w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9858w9859w9860w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9858w9859w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9866w9867w9868w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9866w9867w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9874w9875w9876w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9874w9875w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9882w9883w9884w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9882w9883w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9738w9739w9740w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9738w9739w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9890w9891w9892w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9890w9891w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9898w9899w9900w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9898w9899w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9906w9907w9908w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9906w9907w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9914w9915w9916w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9914w9915w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9922w9923w9924w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9922w9923w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9930w9931w9932w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9930w9931w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9938w9939w9940w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9938w9939w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9946w9947w9948w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9946w9947w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9954w9955w9956w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9954w9955w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9962w9963w9964w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9962w9963w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9746w9747w9748w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9746w9747w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9970w9971w9972w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9970w9971w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9978w9979w9980w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9978w9979w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9754w9755w9756w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9754w9755w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9762w9763w9764w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9762w9763w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9770w9771w9772w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9770w9771w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9778w9779w9780w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9778w9779w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9786w9787w9788w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9786w9787w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9794w9795w9796w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9794w9795w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9802w9803w9804w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_12_w_range9802w9803w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1248w1249w1250w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1248w1249w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1329w1330w1331w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1329w1330w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1337w1338w1339w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1337w1338w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1345w1346w1347w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1345w1346w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1353w1354w1355w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1353w1354w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1361w1362w1363w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1361w1362w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1369w1370w1371w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1369w1370w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1377w1378w1379w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1377w1378w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1385w1386w1387w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1385w1386w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1393w1394w1395w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1393w1394w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1401w1402w1403w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1401w1402w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1257w1258w1259w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1257w1258w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1409w1410w1411w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1409w1410w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1417w1418w1419w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1417w1418w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1425w1426w1427w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1425w1426w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1433w1434w1435w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1433w1434w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1441w1442w1443w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1441w1442w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1449w1450w1451w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1449w1450w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1457w1458w1459w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1457w1458w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1465w1466w1467w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1465w1466w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1473w1474w1475w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1473w1474w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1481w1482w1483w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1481w1482w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1265w1266w1267w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1265w1266w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1489w1490w1491w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1489w1490w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1497w1498w1499w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1497w1498w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1273w1274w1275w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1273w1274w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1281w1282w1283w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1281w1282w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1289w1290w1291w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1289w1290w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1297w1298w1299w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1297w1298w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1305w1306w1307w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1305w1306w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1313w1314w1315w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1313w1314w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1321w1322w1323w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_1_w_range1321w1322w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2044w2045w2046w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2044w2045w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2125w2126w2127w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2125w2126w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2133w2134w2135w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2133w2134w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2141w2142w2143w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2141w2142w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2149w2150w2151w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2149w2150w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2157w2158w2159w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2157w2158w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2165w2166w2167w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2165w2166w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2173w2174w2175w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2173w2174w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2181w2182w2183w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2181w2182w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2189w2190w2191w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2189w2190w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2197w2198w2199w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2197w2198w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2053w2054w2055w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2053w2054w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2205w2206w2207w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2205w2206w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2213w2214w2215w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2213w2214w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2221w2222w2223w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2221w2222w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2229w2230w2231w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2229w2230w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2237w2238w2239w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2237w2238w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2245w2246w2247w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2245w2246w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2253w2254w2255w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2253w2254w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2261w2262w2263w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2261w2262w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2269w2270w2271w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2269w2270w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2277w2278w2279w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2277w2278w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2061w2062w2063w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2061w2062w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2285w2286w2287w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2285w2286w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2293w2294w2295w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2293w2294w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2069w2070w2071w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2069w2070w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2077w2078w2079w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2077w2078w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2085w2086w2087w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2085w2086w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2093w2094w2095w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2093w2094w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2101w2102w2103w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2101w2102w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2109w2110w2111w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2109w2110w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2117w2118w2119w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_2_w_range2117w2118w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2835w2836w2837w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2835w2836w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2916w2917w2918w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2916w2917w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2924w2925w2926w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2924w2925w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2932w2933w2934w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2932w2933w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2940w2941w2942w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2940w2941w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2948w2949w2950w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2948w2949w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2956w2957w2958w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2956w2957w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2964w2965w2966w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2964w2965w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2972w2973w2974w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2972w2973w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2980w2981w2982w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2980w2981w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2988w2989w2990w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2988w2989w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2844w2845w2846w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2844w2845w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2996w2997w2998w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2996w2997w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3004w3005w3006w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3004w3005w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3012w3013w3014w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3012w3013w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3020w3021w3022w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3020w3021w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3028w3029w3030w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3028w3029w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3036w3037w3038w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3036w3037w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3044w3045w3046w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3044w3045w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3052w3053w3054w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3052w3053w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3060w3061w3062w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3060w3061w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3068w3069w3070w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3068w3069w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2852w2853w2854w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2852w2853w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3076w3077w3078w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3076w3077w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3084w3085w3086w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range3084w3085w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2860w2861w2862w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2860w2861w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2868w2869w2870w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2868w2869w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2876w2877w2878w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2876w2877w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2884w2885w2886w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2884w2885w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2892w2893w2894w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2892w2893w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2900w2901w2902w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2900w2901w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2908w2909w2910w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_3_w_range2908w2909w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3621w3622w3623w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3621w3622w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3702w3703w3704w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3702w3703w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3710w3711w3712w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3710w3711w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3718w3719w3720w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3718w3719w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3726w3727w3728w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3726w3727w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3734w3735w3736w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3734w3735w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3742w3743w3744w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3742w3743w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3750w3751w3752w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3750w3751w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3758w3759w3760w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3758w3759w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3766w3767w3768w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3766w3767w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3774w3775w3776w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3774w3775w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3630w3631w3632w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3630w3631w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3782w3783w3784w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3782w3783w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3790w3791w3792w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3790w3791w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3798w3799w3800w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3798w3799w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3806w3807w3808w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3806w3807w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3814w3815w3816w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3814w3815w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3822w3823w3824w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3822w3823w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3830w3831w3832w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3830w3831w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3838w3839w3840w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3838w3839w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3846w3847w3848w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3846w3847w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3854w3855w3856w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3854w3855w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3638w3639w3640w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3638w3639w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3862w3863w3864w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3862w3863w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3870w3871w3872w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3870w3871w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3646w3647w3648w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3646w3647w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3654w3655w3656w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3654w3655w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3662w3663w3664w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3662w3663w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3670w3671w3672w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3670w3671w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3678w3679w3680w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3678w3679w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3686w3687w3688w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3686w3687w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3694w3695w3696w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_4_w_range3694w3695w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4402w4403w4404w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4402w4403w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4483w4484w4485w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4483w4484w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4491w4492w4493w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4491w4492w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4499w4500w4501w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4499w4500w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4507w4508w4509w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4507w4508w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4515w4516w4517w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4515w4516w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4523w4524w4525w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4523w4524w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4531w4532w4533w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4531w4532w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4539w4540w4541w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4539w4540w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4547w4548w4549w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4547w4548w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4555w4556w4557w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4555w4556w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4411w4412w4413w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4411w4412w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4563w4564w4565w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4563w4564w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4571w4572w4573w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4571w4572w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4579w4580w4581w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4579w4580w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4587w4588w4589w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4587w4588w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4595w4596w4597w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4595w4596w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4603w4604w4605w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4603w4604w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4611w4612w4613w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4611w4612w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4619w4620w4621w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4619w4620w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4627w4628w4629w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4627w4628w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4635w4636w4637w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4635w4636w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4419w4420w4421w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4419w4420w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4643w4644w4645w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4643w4644w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4651w4652w4653w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4651w4652w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4427w4428w4429w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4427w4428w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4435w4436w4437w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4435w4436w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4443w4444w4445w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4443w4444w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4451w4452w4453w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4451w4452w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4459w4460w4461w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4459w4460w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4467w4468w4469w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4467w4468w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4475w4476w4477w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_5_w_range4475w4476w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5178w5179w5180w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5178w5179w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5259w5260w5261w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5259w5260w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5267w5268w5269w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5267w5268w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5275w5276w5277w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5275w5276w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5283w5284w5285w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5283w5284w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5291w5292w5293w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5291w5292w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5299w5300w5301w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5299w5300w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5307w5308w5309w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5307w5308w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5315w5316w5317w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5315w5316w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5323w5324w5325w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5323w5324w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5331w5332w5333w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5331w5332w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5187w5188w5189w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5187w5188w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5339w5340w5341w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5339w5340w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5347w5348w5349w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5347w5348w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5355w5356w5357w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5355w5356w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5363w5364w5365w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5363w5364w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5371w5372w5373w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5371w5372w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5379w5380w5381w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5379w5380w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5387w5388w5389w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5387w5388w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5395w5396w5397w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5395w5396w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5403w5404w5405w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5403w5404w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5411w5412w5413w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5411w5412w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5195w5196w5197w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5195w5196w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5419w5420w5421w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5419w5420w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5427w5428w5429w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5427w5428w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5203w5204w5205w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5203w5204w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5211w5212w5213w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5211w5212w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5219w5220w5221w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5219w5220w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5227w5228w5229w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5227w5228w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5235w5236w5237w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5235w5236w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5243w5244w5245w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5243w5244w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5251w5252w5253w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_6_w_range5251w5252w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5949w5950w5951w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5949w5950w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6030w6031w6032w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6030w6031w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6038w6039w6040w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6038w6039w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6046w6047w6048w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6046w6047w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6054w6055w6056w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6054w6055w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6062w6063w6064w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6062w6063w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6070w6071w6072w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6070w6071w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6078w6079w6080w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6078w6079w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6086w6087w6088w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6086w6087w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6094w6095w6096w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6094w6095w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6102w6103w6104w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6102w6103w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5958w5959w5960w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5958w5959w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6110w6111w6112w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6110w6111w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6118w6119w6120w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6118w6119w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6126w6127w6128w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6126w6127w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6134w6135w6136w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6134w6135w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6142w6143w6144w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6142w6143w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6150w6151w6152w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6150w6151w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6158w6159w6160w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6158w6159w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6166w6167w6168w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6166w6167w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6174w6175w6176w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6174w6175w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6182w6183w6184w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6182w6183w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5966w5967w5968w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5966w5967w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6190w6191w6192w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6190w6191w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6198w6199w6200w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6198w6199w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5974w5975w5976w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5974w5975w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5982w5983w5984w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5982w5983w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5990w5991w5992w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5990w5991w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5998w5999w6000w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range5998w5999w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6006w6007w6008w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6006w6007w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6014w6015w6016w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6014w6015w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6022w6023w6024w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_7_w_range6022w6023w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6715w6716w6717w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6715w6716w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6796w6797w6798w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6796w6797w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6804w6805w6806w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6804w6805w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6812w6813w6814w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6812w6813w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6820w6821w6822w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6820w6821w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6828w6829w6830w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6828w6829w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6836w6837w6838w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6836w6837w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6844w6845w6846w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6844w6845w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6852w6853w6854w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6852w6853w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6860w6861w6862w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6860w6861w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6868w6869w6870w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6868w6869w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6724w6725w6726w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6724w6725w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6876w6877w6878w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6876w6877w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6884w6885w6886w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6884w6885w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6892w6893w6894w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6892w6893w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6900w6901w6902w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6900w6901w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6908w6909w6910w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6908w6909w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6916w6917w6918w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6916w6917w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6924w6925w6926w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6924w6925w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6932w6933w6934w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6932w6933w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6940w6941w6942w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6940w6941w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6948w6949w6950w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6948w6949w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6732w6733w6734w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6732w6733w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6956w6957w6958w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6956w6957w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6964w6965w6966w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6964w6965w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6740w6741w6742w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6740w6741w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6748w6749w6750w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6748w6749w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6756w6757w6758w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6756w6757w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6764w6765w6766w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6764w6765w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6772w6773w6774w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6772w6773w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6780w6781w6782w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6780w6781w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6788w6789w6790w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_8_w_range6788w6789w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7476w7477w7478w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7476w7477w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7557w7558w7559w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7557w7558w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7565w7566w7567w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7565w7566w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7573w7574w7575w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7573w7574w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7581w7582w7583w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7581w7582w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7589w7590w7591w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7589w7590w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7597w7598w7599w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7597w7598w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7605w7606w7607w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7605w7606w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7613w7614w7615w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7613w7614w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7621w7622w7623w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7621w7622w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7629w7630w7631w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7629w7630w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7485w7486w7487w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7485w7486w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7637w7638w7639w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7637w7638w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7645w7646w7647w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7645w7646w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7653w7654w7655w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7653w7654w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7661w7662w7663w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7661w7662w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7669w7670w7671w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7669w7670w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7677w7678w7679w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7677w7678w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7685w7686w7687w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7685w7686w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7693w7694w7695w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7693w7694w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7701w7702w7703w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7701w7702w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7709w7710w7711w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7709w7710w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7493w7494w7495w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7493w7494w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7717w7718w7719w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7717w7718w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7725w7726w7727w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7725w7726w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7501w7502w7503w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7501w7502w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7509w7510w7511w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7509w7510w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7517w7518w7519w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7517w7518w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7525w7526w7527w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7525w7526w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7533w7534w7535w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7533w7534w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7541w7542w7543w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7541w7542w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7549w7550w7551w(0) <= wire_ccc_cordic_m_w_lg_w_atannode_9_w_range7549w7550w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	loop31 : FOR i IN 0 TO 31 GENERATE 
		wire_ccc_cordic_m_w_lg_estimate_w10152w(i) <= estimate_w(i) XOR wire_sincosbitff_w_lg_w_q_range9989w9990w(0);
	END GENERATE loop31;
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7214w7470w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7214w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7296w7553w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7296w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7304w7561w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7304w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7312w7569w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7312w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7320w7577w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7320w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7328w7585w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7328w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7336w7593w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7336w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7344w7601w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7344w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7352w7609w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7352w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7360w7617w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7360w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7368w7625w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7368w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7224w7481w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7224w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7376w7633w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7376w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7384w7641w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7384w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7392w7649w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7392w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7400w7657w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7400w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7408w7665w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7408w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7416w7673w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7416w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7424w7681w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7424w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7432w7689w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7432w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7440w7697w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7440w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7448w7705w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7448w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7232w7489w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7232w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7456w7713w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7456w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7464w7721w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7464w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7240w7497w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7240w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7248w7505w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7248w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7256w7513w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7256w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7264w7521w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7264w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7272w7529w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7272w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7280w7537w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7280w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7288w7545w(0) <= wire_ccc_cordic_m_w_x_prenode_10_w_range7288w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range7970w8226w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range7970w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8052w8309w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8052w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8060w8317w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8060w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8068w8325w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8068w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8076w8333w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8076w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8084w8341w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8084w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8092w8349w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8092w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8100w8357w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8100w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8108w8365w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8108w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8116w8373w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8116w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8124w8381w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8124w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range7980w8237w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range7980w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8132w8389w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8132w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8140w8397w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8140w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8148w8405w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8148w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8156w8413w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8156w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8164w8421w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8164w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8172w8429w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8172w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8180w8437w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8180w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8188w8445w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8188w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8196w8453w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8196w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8204w8461w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8204w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range7988w8245w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range7988w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8212w8469w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8212w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8220w8477w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8220w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range7996w8253w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range7996w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8004w8261w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8004w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8012w8269w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8012w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8020w8277w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8020w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8028w8285w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8028w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8036w8293w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8036w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8044w8301w(0) <= wire_ccc_cordic_m_w_x_prenode_11_w_range8044w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8721w8977w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8721w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8803w9060w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8803w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8811w9068w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8811w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8819w9076w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8819w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8827w9084w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8827w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8835w9092w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8835w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8843w9100w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8843w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8851w9108w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8851w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8859w9116w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8859w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8867w9124w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8867w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8875w9132w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8875w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8731w8988w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8731w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8883w9140w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8883w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8891w9148w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8891w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8899w9156w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8899w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8907w9164w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8907w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8915w9172w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8915w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8923w9180w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8923w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8931w9188w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8931w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8939w9196w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8939w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8947w9204w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8947w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8955w9212w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8955w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8739w8996w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8739w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8963w9220w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8963w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8971w9228w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8971w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8747w9004w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8747w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8755w9012w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8755w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8763w9020w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8763w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8771w9028w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8771w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8779w9036w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8779w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8787w9044w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8787w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8795w9052w(0) <= wire_ccc_cordic_m_w_x_prenode_12_w_range8795w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9467w9723w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9467w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9549w9806w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9549w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9557w9814w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9557w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9565w9822w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9565w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9573w9830w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9573w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9581w9838w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9581w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9589w9846w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9589w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9597w9854w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9597w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9605w9862w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9605w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9613w9870w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9613w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9621w9878w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9621w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9477w9734w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9477w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9629w9886w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9629w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9637w9894w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9637w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9645w9902w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9645w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9653w9910w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9653w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9661w9918w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9661w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9669w9926w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9669w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9677w9934w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9677w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9685w9942w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9685w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9693w9950w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9693w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9701w9958w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9701w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9485w9742w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9485w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9709w9966w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9709w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9717w9974w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9717w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9493w9750w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9493w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9501w9758w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9501w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9509w9766w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9509w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9517w9774w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9517w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9525w9782w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9525w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9533w9790w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9533w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9541w9798w(0) <= wire_ccc_cordic_m_w_x_prenode_13_w_range9541w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range986w1242w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range986w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1068w1325w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1068w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1076w1333w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1076w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1084w1341w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1084w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1092w1349w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1092w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1100w1357w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1100w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1108w1365w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1108w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1116w1373w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1116w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1124w1381w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1124w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1132w1389w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1132w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1140w1397w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1140w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range996w1253w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range996w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1148w1405w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1148w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1156w1413w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1156w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1164w1421w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1164w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1172w1429w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1172w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1180w1437w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1180w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1188w1445w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1188w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1196w1453w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1196w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1204w1461w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1204w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1212w1469w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1212w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1220w1477w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1220w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1004w1261w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1004w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1228w1485w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1228w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1236w1493w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1236w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1012w1269w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1012w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1020w1277w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1020w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1028w1285w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1028w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1036w1293w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1036w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1044w1301w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1044w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1052w1309w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1052w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1060w1317w(0) <= wire_ccc_cordic_m_w_x_prenode_2_w_range1060w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1782w2038w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1782w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1864w2121w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1864w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1872w2129w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1872w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1880w2137w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1880w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1888w2145w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1888w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1896w2153w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1896w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1904w2161w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1904w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1912w2169w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1912w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1920w2177w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1920w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1928w2185w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1928w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1936w2193w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1936w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1792w2049w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1792w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1944w2201w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1944w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1952w2209w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1952w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1960w2217w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1960w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1968w2225w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1968w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1976w2233w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1976w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1984w2241w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1984w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1992w2249w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1992w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2000w2257w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2000w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2008w2265w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2008w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2016w2273w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2016w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1800w2057w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1800w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2024w2281w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2024w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2032w2289w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range2032w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1808w2065w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1808w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1816w2073w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1816w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1824w2081w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1824w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1832w2089w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1832w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1840w2097w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1840w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1848w2105w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1848w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1856w2113w(0) <= wire_ccc_cordic_m_w_x_prenode_3_w_range1856w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2573w2829w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2573w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2655w2912w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2655w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2663w2920w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2663w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2671w2928w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2671w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2679w2936w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2679w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2687w2944w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2687w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2695w2952w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2695w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2703w2960w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2703w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2711w2968w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2711w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2719w2976w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2719w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2727w2984w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2727w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2583w2840w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2583w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2735w2992w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2735w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2743w3000w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2743w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2751w3008w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2751w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2759w3016w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2759w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2767w3024w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2767w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2775w3032w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2775w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2783w3040w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2783w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2791w3048w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2791w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2799w3056w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2799w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2807w3064w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2807w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2591w2848w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2591w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2815w3072w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2815w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2823w3080w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2823w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2599w2856w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2599w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2607w2864w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2607w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2615w2872w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2615w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2623w2880w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2623w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2631w2888w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2631w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2639w2896w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2639w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2647w2904w(0) <= wire_ccc_cordic_m_w_x_prenode_4_w_range2647w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3359w3615w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3359w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3441w3698w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3441w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3449w3706w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3449w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3457w3714w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3457w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3465w3722w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3465w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3473w3730w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3473w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3481w3738w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3481w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3489w3746w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3489w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3497w3754w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3497w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3505w3762w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3505w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3513w3770w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3513w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3369w3626w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3369w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3521w3778w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3521w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3529w3786w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3529w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3537w3794w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3537w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3545w3802w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3545w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3553w3810w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3553w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3561w3818w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3561w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3569w3826w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3569w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3577w3834w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3577w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3585w3842w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3585w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3593w3850w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3593w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3377w3634w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3377w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3601w3858w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3601w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3609w3866w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3609w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3385w3642w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3385w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3393w3650w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3393w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3401w3658w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3401w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3409w3666w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3409w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3417w3674w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3417w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3425w3682w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3425w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3433w3690w(0) <= wire_ccc_cordic_m_w_x_prenode_5_w_range3433w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4140w4396w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4140w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4222w4479w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4222w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4230w4487w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4230w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4238w4495w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4238w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4246w4503w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4246w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4254w4511w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4254w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4262w4519w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4262w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4270w4527w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4270w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4278w4535w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4278w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4286w4543w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4286w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4294w4551w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4294w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4150w4407w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4150w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4302w4559w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4302w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4310w4567w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4310w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4318w4575w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4318w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4326w4583w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4326w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4334w4591w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4334w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4342w4599w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4342w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4350w4607w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4350w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4358w4615w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4358w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4366w4623w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4366w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4374w4631w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4374w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4158w4415w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4158w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4382w4639w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4382w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4390w4647w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4390w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4166w4423w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4166w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4174w4431w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4174w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4182w4439w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4182w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4190w4447w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4190w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4198w4455w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4198w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4206w4463w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4206w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4214w4471w(0) <= wire_ccc_cordic_m_w_x_prenode_6_w_range4214w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4916w5172w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range4916w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4998w5255w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range4998w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5006w5263w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5006w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5014w5271w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5014w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5022w5279w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5022w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5030w5287w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5030w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5038w5295w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5038w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5046w5303w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5046w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5054w5311w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5054w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5062w5319w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5062w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5070w5327w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5070w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4926w5183w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range4926w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5078w5335w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5078w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5086w5343w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5086w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5094w5351w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5094w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5102w5359w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5102w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5110w5367w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5110w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5118w5375w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5118w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5126w5383w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5126w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5134w5391w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5134w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5142w5399w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5142w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5150w5407w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5150w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4934w5191w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range4934w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5158w5415w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5158w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5166w5423w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range5166w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4942w5199w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range4942w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4950w5207w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range4950w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4958w5215w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range4958w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4966w5223w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range4966w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4974w5231w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range4974w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4982w5239w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range4982w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4990w5247w(0) <= wire_ccc_cordic_m_w_x_prenode_7_w_range4990w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5687w5943w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5687w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5769w6026w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5769w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5777w6034w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5777w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5785w6042w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5785w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5793w6050w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5793w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5801w6058w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5801w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5809w6066w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5809w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5817w6074w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5817w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5825w6082w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5825w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5833w6090w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5833w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5841w6098w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5841w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5697w5954w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5697w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5849w6106w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5849w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5857w6114w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5857w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5865w6122w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5865w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5873w6130w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5873w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5881w6138w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5881w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5889w6146w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5889w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5897w6154w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5897w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5905w6162w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5905w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5913w6170w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5913w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5921w6178w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5921w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5705w5962w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5705w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5929w6186w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5929w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5937w6194w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5937w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5713w5970w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5713w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5721w5978w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5721w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5729w5986w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5729w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5737w5994w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5737w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5745w6002w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5745w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5753w6010w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5753w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5761w6018w(0) <= wire_ccc_cordic_m_w_x_prenode_8_w_range5761w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6453w6709w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6453w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6535w6792w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6535w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6543w6800w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6543w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6551w6808w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6551w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6559w6816w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6559w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6567w6824w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6567w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6575w6832w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6575w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6583w6840w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6583w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6591w6848w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6591w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6599w6856w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6599w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6607w6864w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6607w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6463w6720w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6463w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6615w6872w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6615w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6623w6880w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6623w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6631w6888w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6631w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6639w6896w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6639w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6647w6904w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6647w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6655w6912w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6655w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6663w6920w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6663w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6671w6928w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6671w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6679w6936w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6679w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6687w6944w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6687w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6471w6728w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6471w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6695w6952w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6695w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6703w6960w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6703w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6479w6736w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6479w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6487w6744w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6487w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6495w6752w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6495w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6503w6760w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6503w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6511w6768w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6511w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6519w6776w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6519w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6527w6784w(0) <= wire_ccc_cordic_m_w_x_prenode_9_w_range6527w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7219w7473w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7219w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7300w7555w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7300w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7308w7563w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7308w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7316w7571w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7316w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7324w7579w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7324w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7332w7587w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7332w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7340w7595w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7340w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7348w7603w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7348w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7356w7611w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7356w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7364w7619w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7364w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7372w7627w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7372w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7228w7483w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7228w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7380w7635w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7380w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7388w7643w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7388w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7396w7651w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7396w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7404w7659w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7404w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7412w7667w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7412w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7420w7675w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7420w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7428w7683w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7428w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7436w7691w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7436w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7444w7699w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7444w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7452w7707w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7452w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7236w7491w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7236w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7460w7715w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7460w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7468w7723w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7468w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7244w7499w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7244w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7252w7507w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7252w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7260w7515w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7260w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7268w7523w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7268w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7276w7531w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7276w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7284w7539w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7284w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7292w7547w(0) <= wire_ccc_cordic_m_w_y_prenode_10_w_range7292w(0) XOR wire_z_pipeff_9_w_q_range7469w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range7975w8229w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range7975w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8056w8311w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8056w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8064w8319w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8064w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8072w8327w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8072w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8080w8335w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8080w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8088w8343w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8088w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8096w8351w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8096w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8104w8359w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8104w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8112w8367w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8112w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8120w8375w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8120w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8128w8383w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8128w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range7984w8239w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range7984w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8136w8391w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8136w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8144w8399w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8144w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8152w8407w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8152w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8160w8415w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8160w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8168w8423w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8168w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8176w8431w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8176w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8184w8439w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8184w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8192w8447w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8192w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8200w8455w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8200w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8208w8463w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8208w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range7992w8247w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range7992w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8216w8471w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8216w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8224w8479w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8224w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8000w8255w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8000w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8008w8263w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8008w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8016w8271w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8016w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8024w8279w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8024w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8032w8287w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8032w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8040w8295w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8040w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8048w8303w(0) <= wire_ccc_cordic_m_w_y_prenode_11_w_range8048w(0) XOR wire_z_pipeff_10_w_q_range8225w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8726w8980w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8726w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8807w9062w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8807w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8815w9070w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8815w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8823w9078w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8823w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8831w9086w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8831w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8839w9094w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8839w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8847w9102w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8847w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8855w9110w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8855w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8863w9118w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8863w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8871w9126w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8871w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8879w9134w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8879w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8735w8990w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8735w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8887w9142w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8887w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8895w9150w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8895w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8903w9158w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8903w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8911w9166w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8911w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8919w9174w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8919w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8927w9182w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8927w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8935w9190w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8935w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8943w9198w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8943w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8951w9206w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8951w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8959w9214w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8959w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8743w8998w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8743w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8967w9222w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8967w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8975w9230w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8975w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8751w9006w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8751w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8759w9014w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8759w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8767w9022w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8767w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8775w9030w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8775w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8783w9038w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8783w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8791w9046w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8791w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8799w9054w(0) <= wire_ccc_cordic_m_w_y_prenode_12_w_range8799w(0) XOR wire_z_pipeff_11_w_q_range8976w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9472w9726w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9472w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9553w9808w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9553w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9561w9816w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9561w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9569w9824w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9569w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9577w9832w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9577w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9585w9840w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9585w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9593w9848w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9593w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9601w9856w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9601w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9609w9864w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9609w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9617w9872w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9617w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9625w9880w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9625w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9481w9736w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9481w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9633w9888w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9633w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9641w9896w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9641w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9649w9904w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9649w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9657w9912w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9657w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9665w9920w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9665w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9673w9928w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9673w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9681w9936w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9681w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9689w9944w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9689w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9697w9952w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9697w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9705w9960w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9705w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9489w9744w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9489w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9713w9968w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9713w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9721w9976w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9721w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9497w9752w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9497w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9505w9760w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9505w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9513w9768w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9513w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9521w9776w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9521w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9529w9784w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9529w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9537w9792w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9537w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9545w9800w(0) <= wire_ccc_cordic_m_w_y_prenode_13_w_range9545w(0) XOR wire_z_pipeff_12_w_q_range9722w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range991w1245w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range991w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1072w1327w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1072w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1080w1335w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1080w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1088w1343w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1088w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1096w1351w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1096w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1104w1359w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1104w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1112w1367w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1112w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1120w1375w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1120w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1128w1383w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1128w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1136w1391w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1136w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1144w1399w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1144w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1000w1255w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1000w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1152w1407w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1152w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1160w1415w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1160w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1168w1423w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1168w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1176w1431w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1176w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1184w1439w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1184w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1192w1447w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1192w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1200w1455w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1200w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1208w1463w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1208w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1216w1471w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1216w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1224w1479w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1224w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1008w1263w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1008w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1232w1487w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1232w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1240w1495w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1240w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1016w1271w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1016w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1024w1279w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1024w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1032w1287w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1032w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1040w1295w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1040w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1048w1303w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1048w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1056w1311w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1056w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1064w1319w(0) <= wire_ccc_cordic_m_w_y_prenode_2_w_range1064w(0) XOR wire_z_pipeff_1_w_q_range1241w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1787w2041w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1787w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1868w2123w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1868w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1876w2131w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1876w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1884w2139w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1884w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1892w2147w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1892w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1900w2155w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1900w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1908w2163w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1908w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1916w2171w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1916w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1924w2179w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1924w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1932w2187w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1932w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1940w2195w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1940w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1796w2051w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1796w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1948w2203w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1948w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1956w2211w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1956w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1964w2219w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1964w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1972w2227w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1972w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1980w2235w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1980w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1988w2243w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1988w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1996w2251w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1996w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2004w2259w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2004w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2012w2267w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2012w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2020w2275w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2020w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1804w2059w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1804w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2028w2283w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2028w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2036w2291w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range2036w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1812w2067w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1812w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1820w2075w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1820w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1828w2083w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1828w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1836w2091w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1836w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1844w2099w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1844w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1852w2107w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1852w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1860w2115w(0) <= wire_ccc_cordic_m_w_y_prenode_3_w_range1860w(0) XOR wire_z_pipeff_2_w_q_range2037w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2578w2832w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2578w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2659w2914w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2659w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2667w2922w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2667w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2675w2930w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2675w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2683w2938w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2683w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2691w2946w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2691w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2699w2954w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2699w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2707w2962w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2707w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2715w2970w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2715w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2723w2978w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2723w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2731w2986w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2731w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2587w2842w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2587w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2739w2994w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2739w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2747w3002w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2747w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2755w3010w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2755w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2763w3018w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2763w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2771w3026w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2771w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2779w3034w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2779w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2787w3042w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2787w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2795w3050w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2795w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2803w3058w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2803w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2811w3066w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2811w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2595w2850w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2595w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2819w3074w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2819w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2827w3082w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2827w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2603w2858w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2603w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2611w2866w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2611w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2619w2874w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2619w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2627w2882w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2627w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2635w2890w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2635w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2643w2898w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2643w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2651w2906w(0) <= wire_ccc_cordic_m_w_y_prenode_4_w_range2651w(0) XOR wire_z_pipeff_3_w_q_range2828w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3364w3618w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3364w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3445w3700w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3445w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3453w3708w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3453w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3461w3716w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3461w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3469w3724w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3469w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3477w3732w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3477w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3485w3740w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3485w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3493w3748w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3493w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3501w3756w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3501w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3509w3764w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3509w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3517w3772w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3517w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3373w3628w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3373w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3525w3780w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3525w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3533w3788w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3533w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3541w3796w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3541w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3549w3804w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3549w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3557w3812w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3557w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3565w3820w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3565w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3573w3828w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3573w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3581w3836w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3581w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3589w3844w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3589w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3597w3852w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3597w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3381w3636w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3381w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3605w3860w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3605w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3613w3868w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3613w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3389w3644w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3389w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3397w3652w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3397w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3405w3660w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3405w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3413w3668w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3413w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3421w3676w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3421w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3429w3684w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3429w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3437w3692w(0) <= wire_ccc_cordic_m_w_y_prenode_5_w_range3437w(0) XOR wire_z_pipeff_4_w_q_range3614w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4145w4399w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4145w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4226w4481w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4226w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4234w4489w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4234w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4242w4497w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4242w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4250w4505w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4250w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4258w4513w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4258w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4266w4521w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4266w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4274w4529w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4274w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4282w4537w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4282w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4290w4545w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4290w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4298w4553w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4298w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4154w4409w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4154w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4306w4561w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4306w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4314w4569w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4314w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4322w4577w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4322w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4330w4585w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4330w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4338w4593w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4338w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4346w4601w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4346w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4354w4609w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4354w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4362w4617w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4362w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4370w4625w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4370w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4378w4633w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4378w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4162w4417w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4162w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4386w4641w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4386w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4394w4649w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4394w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4170w4425w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4170w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4178w4433w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4178w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4186w4441w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4186w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4194w4449w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4194w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4202w4457w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4202w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4210w4465w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4210w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4218w4473w(0) <= wire_ccc_cordic_m_w_y_prenode_6_w_range4218w(0) XOR wire_z_pipeff_5_w_q_range4395w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4921w5175w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range4921w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5002w5257w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5002w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5010w5265w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5010w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5018w5273w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5018w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5026w5281w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5026w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5034w5289w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5034w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5042w5297w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5042w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5050w5305w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5050w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5058w5313w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5058w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5066w5321w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5066w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5074w5329w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5074w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4930w5185w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range4930w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5082w5337w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5082w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5090w5345w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5090w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5098w5353w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5098w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5106w5361w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5106w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5114w5369w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5114w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5122w5377w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5122w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5130w5385w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5130w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5138w5393w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5138w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5146w5401w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5146w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5154w5409w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5154w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4938w5193w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range4938w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5162w5417w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5162w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5170w5425w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range5170w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4946w5201w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range4946w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4954w5209w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range4954w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4962w5217w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range4962w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4970w5225w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range4970w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4978w5233w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range4978w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4986w5241w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range4986w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4994w5249w(0) <= wire_ccc_cordic_m_w_y_prenode_7_w_range4994w(0) XOR wire_z_pipeff_6_w_q_range5171w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5692w5946w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5692w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5773w6028w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5773w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5781w6036w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5781w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5789w6044w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5789w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5797w6052w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5797w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5805w6060w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5805w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5813w6068w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5813w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5821w6076w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5821w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5829w6084w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5829w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5837w6092w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5837w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5845w6100w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5845w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5701w5956w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5701w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5853w6108w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5853w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5861w6116w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5861w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5869w6124w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5869w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5877w6132w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5877w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5885w6140w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5885w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5893w6148w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5893w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5901w6156w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5901w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5909w6164w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5909w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5917w6172w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5917w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5925w6180w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5925w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5709w5964w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5709w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5933w6188w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5933w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5941w6196w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5941w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5717w5972w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5717w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5725w5980w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5725w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5733w5988w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5733w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5741w5996w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5741w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5749w6004w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5749w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5757w6012w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5757w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5765w6020w(0) <= wire_ccc_cordic_m_w_y_prenode_8_w_range5765w(0) XOR wire_z_pipeff_7_w_q_range5942w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6458w6712w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6458w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6539w6794w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6539w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6547w6802w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6547w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6555w6810w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6555w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6563w6818w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6563w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6571w6826w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6571w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6579w6834w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6579w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6587w6842w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6587w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6595w6850w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6595w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6603w6858w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6603w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6611w6866w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6611w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6467w6722w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6467w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6619w6874w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6619w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6627w6882w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6627w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6635w6890w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6635w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6643w6898w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6643w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6651w6906w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6651w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6659w6914w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6659w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6667w6922w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6667w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6675w6930w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6675w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6683w6938w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6683w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6691w6946w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6691w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6475w6730w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6475w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6699w6954w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6699w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6707w6962w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6707w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6483w6738w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6483w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6491w6746w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6491w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6499w6754w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6499w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6507w6762w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6507w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6515w6770w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6515w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6523w6778w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6523w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6531w6786w(0) <= wire_ccc_cordic_m_w_y_prenode_9_w_range6531w(0) XOR wire_z_pipeff_8_w_q_range6708w(0);
	atannode_0_w <= wire_cata_0_cordic_atan_arctan;
	atannode_10_w <= wire_cata_10_cordic_atan_arctan;
	atannode_11_w <= wire_cata_11_cordic_atan_arctan;
	atannode_12_w <= wire_cata_12_cordic_atan_arctan;
	atannode_1_w <= wire_cata_1_cordic_atan_arctan;
	atannode_2_w <= wire_cata_2_cordic_atan_arctan;
	atannode_3_w <= wire_cata_3_cordic_atan_arctan;
	atannode_4_w <= wire_cata_4_cordic_atan_arctan;
	atannode_5_w <= wire_cata_5_cordic_atan_arctan;
	atannode_6_w <= wire_cata_6_cordic_atan_arctan;
	atannode_7_w <= wire_cata_7_cordic_atan_arctan;
	atannode_8_w <= wire_cata_8_cordic_atan_arctan;
	atannode_9_w <= wire_cata_9_cordic_atan_arctan;
	delay_input_w <= (wire_x_pipeff_13_w_lg_q9987w OR wire_y_pipeff_13_w_lg_q9986w);
	delay_pipe_w <= cdaff_2;
	estimate_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10138w10149w10150w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10133w10146w10147w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10128w10143w10144w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10123w10140w10141w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10118w10135w10136w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10113w10130w10131w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10108w10125w10126w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10103w10120w10121w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10098w10115w10116w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10093w10110w10111w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10088w10105w10106w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10083w10100w10101w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10078w10095w10096w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10073w10090w10091w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10068w10085w10086w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10063w10080w10081w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10058w10075w10076w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10053w10070w10071w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10048w10065w10066w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10043w10060w10061w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10038w10055w10056w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10033w10050w10051w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10028w10045w10046w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10023w10040w10041w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10018w10035w10036w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10013w10030w10031w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10007w10025w10026w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10001w10020w10021w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range9993w10015w10016w
 & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10009w10010w10011w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range10003w10004w10005w & wire_ccc_cordic_m_w_lg_w_lg_w_pre_estimate_w_range9996w9997w9998w);
	indexpointnum_w <= "0001";
	multiplier_input_w <= (wire_x_pipeff_13_w_lg_q9984w OR wire_y_pipeff_13_w_lg_q9983w);
	multipliernode_w <= wire_cmx_result;
	post_estimate_w <= wire_ccc_cordic_m_w_lg_estimate_w10152w;
	pre_estimate_w <= multipliernode_w(61 DOWNTO 30);
	radians_load_node_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_radians_range440w443w444w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range435w438w439w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range430w433w434w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range425w428w429w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range420w423w424w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range415w418w419w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range410w413w414w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range405w408w409w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range400w403w404w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range395w398w399w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range390w393w394w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range385w388w389w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range380w383w384w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range375w378w379w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range370w373w374w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range365w368w369w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range360w363w364w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range355w358w359w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range350w353w354w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range345w348w349w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range340w343w344w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range335w338w339w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range330w333w334w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range325w328w329w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range320w323w324w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range315w318w319w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range310w313w314w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range305w308w309w & wire_ccc_cordic_m_w_lg_w_lg_w_radians_range300w303w304w & wire_ccc_cordic_m_w_lg_w_radians_range297w299w & wire_ccc_cordic_m_w_lg_w_radians_range294w296w & wire_ccc_cordic_m_w_lg_w_radians_range289w292w);
	sincos <= sincosff;
	startindex_w <= wire_ccc_cordic_m_w_lg_indexpointnum_w288w;
	x_pipenode_10_w <= wire_x_pipenode_10_add_result;
	x_pipenode_11_w <= wire_x_pipenode_11_add_result;
	x_pipenode_12_w <= wire_x_pipenode_12_add_result;
	x_pipenode_13_w <= wire_x_pipenode_13_add_result;
	x_pipenode_2_w <= wire_x_pipenode_2_add_result;
	x_pipenode_3_w <= wire_x_pipenode_3_add_result;
	x_pipenode_4_w <= wire_x_pipenode_4_add_result;
	x_pipenode_5_w <= wire_x_pipenode_5_add_result;
	x_pipenode_6_w <= wire_x_pipenode_6_add_result;
	x_pipenode_7_w <= wire_x_pipenode_7_add_result;
	x_pipenode_8_w <= wire_x_pipenode_8_add_result;
	x_pipenode_9_w <= wire_x_pipenode_9_add_result;
	x_prenode_10_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6989w7462w7463w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6987w7454w7455w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6985w7446w7447w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6983w7438w7439w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6981w7430w7431w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6979w7422w7423w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6977w7414w7415w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6975w7406w7407w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range6970w7398w7399w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7148w7390w7391w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7144w7382w7383w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7138w7374w7375w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7132w7366w7367w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7126w7358w7359w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7120w7350w7351w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7114w7342w7343w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7108w7334w7335w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7102w7326w7327w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7096w7318w7319w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7090w7310w7311w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7084w7302w7303w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7078w7294w7295w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7072w7286w7287w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7066w7278w7279w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7060w7270w7271w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7054w7262w7263w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7048w7254w7255w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7042w7246w7247w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7036w7238w7239w
 & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7030w7230w7231w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7024w7222w7223w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_10_w_range7019w7212w7213w);
	x_prenode_11_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7752w8218w8219w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7750w8210w8211w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7748w8202w8203w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7746w8194w8195w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7744w8186w8187w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7742w8178w8179w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7740w8170w8171w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7738w8162w8163w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7736w8154w8155w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7731w8146w8147w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7907w8138w8139w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7903w8130w8131w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7897w8122w8123w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7891w8114w8115w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7885w8106w8107w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7879w8098w8099w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7873w8090w8091w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7867w8082w8083w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7861w8074w8075w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7855w8066w8067w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7849w8058w8059w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7843w8050w8051w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7837w8042w8043w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7831w8034w8035w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7825w8026w8027w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7819w8018w8019w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7813w8010w8011w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7807w8002w8003w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7801w7994w7995w
 & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7795w7986w7987w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7789w7978w7979w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_11_w_range7784w7968w7969w);
	x_prenode_12_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8510w8969w8970w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8508w8961w8962w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8506w8953w8954w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8504w8945w8946w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8502w8937w8938w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8500w8929w8930w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8498w8921w8922w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8496w8913w8914w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8494w8905w8906w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8492w8897w8898w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8487w8889w8890w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8661w8881w8882w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8657w8873w8874w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8651w8865w8866w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8645w8857w8858w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8639w8849w8850w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8633w8841w8842w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8627w8833w8834w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8621w8825w8826w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8615w8817w8818w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8609w8809w8810w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8603w8801w8802w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8597w8793w8794w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8591w8785w8786w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8585w8777w8778w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8579w8769w8770w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8573w8761w8762w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8567w8753w8754w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8561w8745w8746w
 & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8555w8737w8738w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8549w8729w8730w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_12_w_range8544w8719w8720w);
	x_prenode_13_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9263w9715w9716w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9261w9707w9708w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9259w9699w9700w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9257w9691w9692w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9255w9683w9684w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9253w9675w9676w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9251w9667w9668w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9249w9659w9660w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9247w9651w9652w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9245w9643w9644w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9243w9635w9636w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9238w9627w9628w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9410w9619w9620w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9406w9611w9612w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9400w9603w9604w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9394w9595w9596w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9388w9587w9588w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9382w9579w9580w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9376w9571w9572w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9370w9563w9564w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9364w9555w9556w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9358w9547w9548w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9352w9539w9540w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9346w9531w9532w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9340w9523w9524w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9334w9515w9516w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9328w9507w9508w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9322w9499w9500w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9316w9491w9492w
 & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9310w9483w9484w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9304w9475w9476w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_13_w_range9299w9465w9466w);
	x_prenode_2_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range702w1234w1235w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range896w1226w1227w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range892w1218w1219w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range886w1210w1211w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range880w1202w1203w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range874w1194w1195w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range868w1186w1187w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range862w1178w1179w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range856w1170w1171w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range850w1162w1163w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range844w1154w1155w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range838w1146w1147w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range832w1138w1139w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range826w1130w1131w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range820w1122w1123w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range814w1114w1115w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range808w1106w1107w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range802w1098w1099w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range796w1090w1091w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range790w1082w1083w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range784w1074w1075w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range778w1066w1067w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range772w1058w1059w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range766w1050w1051w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range760w1042w1043w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range754w1034w1035w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range748w1026w1027w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range742w1018w1019w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range736w1010w1011w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range730w1002w1003w
 & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range724w994w995w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_2_w_range719w984w985w);
	x_prenode_3_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1508w2030w2031w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1503w2022w2023w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1695w2014w2015w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1691w2006w2007w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1685w1998w1999w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1679w1990w1991w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1673w1982w1983w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1667w1974w1975w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1661w1966w1967w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1655w1958w1959w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1649w1950w1951w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1643w1942w1943w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1637w1934w1935w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1631w1926w1927w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1625w1918w1919w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1619w1910w1911w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1613w1902w1903w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1607w1894w1895w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1601w1886w1887w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1595w1878w1879w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1589w1870w1871w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1583w1862w1863w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1577w1854w1855w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1571w1846w1847w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1565w1838w1839w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1559w1830w1831w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1553w1822w1823w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1547w1814w1815w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1541w1806w1807w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1535w1798w1799w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1529w1790w1791w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_3_w_range1524w1780w1781w);
	x_prenode_4_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2306w2821w2822w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2304w2813w2814w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2299w2805w2806w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2489w2797w2798w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2485w2789w2790w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2479w2781w2782w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2473w2773w2774w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2467w2765w2766w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2461w2757w2758w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2455w2749w2750w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2449w2741w2742w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2443w2733w2734w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2437w2725w2726w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2431w2717w2718w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2425w2709w2710w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2419w2701w2702w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2413w2693w2694w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2407w2685w2686w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2401w2677w2678w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2395w2669w2670w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2389w2661w2662w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2383w2653w2654w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2377w2645w2646w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2371w2637w2638w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2365w2629w2630w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2359w2621w2622w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2353w2613w2614w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2347w2605w2606w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2341w2597w2598w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2335w2589w2590w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2329w2581w2582w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_4_w_range2324w2571w2572w);
	x_prenode_5_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3099w3607w3608w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3097w3599w3600w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3095w3591w3592w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3090w3583w3584w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3278w3575w3576w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3274w3567w3568w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3268w3559w3560w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3262w3551w3552w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3256w3543w3544w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3250w3535w3536w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3244w3527w3528w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3238w3519w3520w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3232w3511w3512w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3226w3503w3504w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3220w3495w3496w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3214w3487w3488w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3208w3479w3480w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3202w3471w3472w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3196w3463w3464w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3190w3455w3456w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3184w3447w3448w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3178w3439w3440w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3172w3431w3432w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3166w3423w3424w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3160w3415w3416w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3154w3407w3408w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3148w3399w3400w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3142w3391w3392w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3136w3383w3384w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3130w3375w3376w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3124w3367w3368w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_5_w_range3119w3357w3358w);
	x_prenode_6_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3887w4388w4389w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3885w4380w4381w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3883w4372w4373w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3881w4364w4365w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3876w4356w4357w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4062w4348w4349w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4058w4340w4341w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4052w4332w4333w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4046w4324w4325w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4040w4316w4317w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4034w4308w4309w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4028w4300w4301w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4022w4292w4293w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4016w4284w4285w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4010w4276w4277w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range4004w4268w4269w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3998w4260w4261w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3992w4252w4253w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3986w4244w4245w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3980w4236w4237w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3974w4228w4229w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3968w4220w4221w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3962w4212w4213w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3956w4204w4205w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3950w4196w4197w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3944w4188w4189w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3938w4180w4181w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3932w4172w4173w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3926w4164w4165w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3920w4156w4157w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3914w4148w4149w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_6_w_range3909w4138w4139w);
	x_prenode_7_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4670w5164w5165w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4668w5156w5157w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4666w5148w5149w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4664w5140w5141w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4662w5132w5133w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4657w5124w5125w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4841w5116w5117w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4837w5108w5109w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4831w5100w5101w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4825w5092w5093w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4819w5084w5085w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4813w5076w5077w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4807w5068w5069w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4801w5060w5061w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4795w5052w5053w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4789w5044w5045w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4783w5036w5037w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4777w5028w5029w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4771w5020w5021w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4765w5012w5013w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4759w5004w5005w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4753w4996w4997w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4747w4988w4989w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4741w4980w4981w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4735w4972w4973w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4729w4964w4965w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4723w4956w4957w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4717w4948w4949w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4711w4940w4941w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4705w4932w4933w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4699w4924w4925w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_7_w_range4694w4914w4915w);
	x_prenode_8_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5448w5935w5936w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5446w5927w5928w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5444w5919w5920w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5442w5911w5912w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5440w5903w5904w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5438w5895w5896w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5433w5887w5888w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5615w5879w5880w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5611w5871w5872w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5605w5863w5864w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5599w5855w5856w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5593w5847w5848w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5587w5839w5840w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5581w5831w5832w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5575w5823w5824w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5569w5815w5816w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5563w5807w5808w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5557w5799w5800w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5551w5791w5792w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5545w5783w5784w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5539w5775w5776w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5533w5767w5768w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5527w5759w5760w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5521w5751w5752w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5515w5743w5744w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5509w5735w5736w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5503w5727w5728w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5497w5719w5720w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5491w5711w5712w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5485w5703w5704w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5479w5695w5696w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_8_w_range5474w5685w5686w);
	x_prenode_9_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6221w6701w6702w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6219w6693w6694w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6217w6685w6686w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6215w6677w6678w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6213w6669w6670w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6211w6661w6662w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6209w6653w6654w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6204w6645w6646w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6384w6637w6638w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6380w6629w6630w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6374w6621w6622w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6368w6613w6614w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6362w6605w6606w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6356w6597w6598w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6350w6589w6590w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6344w6581w6582w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6338w6573w6574w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6332w6565w6566w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6326w6557w6558w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6320w6549w6550w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6314w6541w6542w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6308w6533w6534w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6302w6525w6526w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6296w6517w6518w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6290w6509w6510w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6284w6501w6502w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6278w6493w6494w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6272w6485w6486w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6266w6477w6478w 
& wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6260w6469w6470w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6254w6461w6462w & wire_ccc_cordic_m_w_lg_w_lg_w_x_prenodeone_9_w_range6249w6451w6452w);
	x_prenodeone_10_w <= ( wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range7142w7143w & wire_y_pipeff_9_w_lg_w_q_range7136w7137w & wire_y_pipeff_9_w_lg_w_q_range7130w7131w & wire_y_pipeff_9_w_lg_w_q_range7124w7125w & wire_y_pipeff_9_w_lg_w_q_range7118w7119w & wire_y_pipeff_9_w_lg_w_q_range7112w7113w & wire_y_pipeff_9_w_lg_w_q_range7106w7107w & wire_y_pipeff_9_w_lg_w_q_range7100w7101w & wire_y_pipeff_9_w_lg_w_q_range7094w7095w & wire_y_pipeff_9_w_lg_w_q_range7088w7089w & wire_y_pipeff_9_w_lg_w_q_range7082w7083w & wire_y_pipeff_9_w_lg_w_q_range7076w7077w & wire_y_pipeff_9_w_lg_w_q_range7070w7071w & wire_y_pipeff_9_w_lg_w_q_range7064w7065w & wire_y_pipeff_9_w_lg_w_q_range7058w7059w & wire_y_pipeff_9_w_lg_w_q_range7052w7053w & wire_y_pipeff_9_w_lg_w_q_range7046w7047w & wire_y_pipeff_9_w_lg_w_q_range7040w7041w & wire_y_pipeff_9_w_lg_w_q_range7034w7035w & wire_y_pipeff_9_w_lg_w_q_range7028w7029w & wire_y_pipeff_9_w_lg_w_q_range7022w7023w & wire_y_pipeff_9_w_lg_w_q_range7017w7018w);
	x_prenodeone_11_w <= ( wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7901w7902w & wire_y_pipeff_10_w_lg_w_q_range7895w7896w & wire_y_pipeff_10_w_lg_w_q_range7889w7890w & wire_y_pipeff_10_w_lg_w_q_range7883w7884w & wire_y_pipeff_10_w_lg_w_q_range7877w7878w & wire_y_pipeff_10_w_lg_w_q_range7871w7872w & wire_y_pipeff_10_w_lg_w_q_range7865w7866w & wire_y_pipeff_10_w_lg_w_q_range7859w7860w & wire_y_pipeff_10_w_lg_w_q_range7853w7854w & wire_y_pipeff_10_w_lg_w_q_range7847w7848w & wire_y_pipeff_10_w_lg_w_q_range7841w7842w & wire_y_pipeff_10_w_lg_w_q_range7835w7836w & wire_y_pipeff_10_w_lg_w_q_range7829w7830w & wire_y_pipeff_10_w_lg_w_q_range7823w7824w & wire_y_pipeff_10_w_lg_w_q_range7817w7818w & wire_y_pipeff_10_w_lg_w_q_range7811w7812w & wire_y_pipeff_10_w_lg_w_q_range7805w7806w & wire_y_pipeff_10_w_lg_w_q_range7799w7800w & wire_y_pipeff_10_w_lg_w_q_range7793w7794w & wire_y_pipeff_10_w_lg_w_q_range7787w7788w & wire_y_pipeff_10_w_lg_w_q_range7782w7783w);
	x_prenodeone_12_w <= ( wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8655w8656w & wire_y_pipeff_11_w_lg_w_q_range8649w8650w & wire_y_pipeff_11_w_lg_w_q_range8643w8644w & wire_y_pipeff_11_w_lg_w_q_range8637w8638w & wire_y_pipeff_11_w_lg_w_q_range8631w8632w & wire_y_pipeff_11_w_lg_w_q_range8625w8626w & wire_y_pipeff_11_w_lg_w_q_range8619w8620w & wire_y_pipeff_11_w_lg_w_q_range8613w8614w & wire_y_pipeff_11_w_lg_w_q_range8607w8608w & wire_y_pipeff_11_w_lg_w_q_range8601w8602w & wire_y_pipeff_11_w_lg_w_q_range8595w8596w & wire_y_pipeff_11_w_lg_w_q_range8589w8590w & wire_y_pipeff_11_w_lg_w_q_range8583w8584w & wire_y_pipeff_11_w_lg_w_q_range8577w8578w & wire_y_pipeff_11_w_lg_w_q_range8571w8572w & wire_y_pipeff_11_w_lg_w_q_range8565w8566w & wire_y_pipeff_11_w_lg_w_q_range8559w8560w & wire_y_pipeff_11_w_lg_w_q_range8553w8554w & wire_y_pipeff_11_w_lg_w_q_range8547w8548w & wire_y_pipeff_11_w_lg_w_q_range8542w8543w);
	x_prenodeone_13_w <= ( wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9404w9405w & wire_y_pipeff_12_w_lg_w_q_range9398w9399w & wire_y_pipeff_12_w_lg_w_q_range9392w9393w & wire_y_pipeff_12_w_lg_w_q_range9386w9387w & wire_y_pipeff_12_w_lg_w_q_range9380w9381w & wire_y_pipeff_12_w_lg_w_q_range9374w9375w & wire_y_pipeff_12_w_lg_w_q_range9368w9369w & wire_y_pipeff_12_w_lg_w_q_range9362w9363w & wire_y_pipeff_12_w_lg_w_q_range9356w9357w & wire_y_pipeff_12_w_lg_w_q_range9350w9351w & wire_y_pipeff_12_w_lg_w_q_range9344w9345w & wire_y_pipeff_12_w_lg_w_q_range9338w9339w & wire_y_pipeff_12_w_lg_w_q_range9332w9333w & wire_y_pipeff_12_w_lg_w_q_range9326w9327w & wire_y_pipeff_12_w_lg_w_q_range9320w9321w & wire_y_pipeff_12_w_lg_w_q_range9314w9315w & wire_y_pipeff_12_w_lg_w_q_range9308w9309w & wire_y_pipeff_12_w_lg_w_q_range9302w9303w & wire_y_pipeff_12_w_lg_w_q_range9297w9298w);
	x_prenodeone_2_w <= ( wire_y_pipeff_1_w_lg_w_q_range700w701w & wire_y_pipeff_1_w_lg_w_q_range700w701w & wire_y_pipeff_1_w_lg_w_q_range890w891w & wire_y_pipeff_1_w_lg_w_q_range884w885w & wire_y_pipeff_1_w_lg_w_q_range878w879w & wire_y_pipeff_1_w_lg_w_q_range872w873w & wire_y_pipeff_1_w_lg_w_q_range866w867w & wire_y_pipeff_1_w_lg_w_q_range860w861w & wire_y_pipeff_1_w_lg_w_q_range854w855w & wire_y_pipeff_1_w_lg_w_q_range848w849w & wire_y_pipeff_1_w_lg_w_q_range842w843w & wire_y_pipeff_1_w_lg_w_q_range836w837w & wire_y_pipeff_1_w_lg_w_q_range830w831w & wire_y_pipeff_1_w_lg_w_q_range824w825w & wire_y_pipeff_1_w_lg_w_q_range818w819w & wire_y_pipeff_1_w_lg_w_q_range812w813w & wire_y_pipeff_1_w_lg_w_q_range806w807w & wire_y_pipeff_1_w_lg_w_q_range800w801w & wire_y_pipeff_1_w_lg_w_q_range794w795w & wire_y_pipeff_1_w_lg_w_q_range788w789w & wire_y_pipeff_1_w_lg_w_q_range782w783w & wire_y_pipeff_1_w_lg_w_q_range776w777w & wire_y_pipeff_1_w_lg_w_q_range770w771w & wire_y_pipeff_1_w_lg_w_q_range764w765w & wire_y_pipeff_1_w_lg_w_q_range758w759w & wire_y_pipeff_1_w_lg_w_q_range752w753w & wire_y_pipeff_1_w_lg_w_q_range746w747w & wire_y_pipeff_1_w_lg_w_q_range740w741w & wire_y_pipeff_1_w_lg_w_q_range734w735w & wire_y_pipeff_1_w_lg_w_q_range728w729w & wire_y_pipeff_1_w_lg_w_q_range722w723w & wire_y_pipeff_1_w_lg_w_q_range717w718w);
	x_prenodeone_3_w <= ( wire_y_pipeff_2_w_lg_w_q_range1501w1502w & wire_y_pipeff_2_w_lg_w_q_range1501w1502w & wire_y_pipeff_2_w_lg_w_q_range1501w1502w & wire_y_pipeff_2_w_lg_w_q_range1689w1690w & wire_y_pipeff_2_w_lg_w_q_range1683w1684w & wire_y_pipeff_2_w_lg_w_q_range1677w1678w & wire_y_pipeff_2_w_lg_w_q_range1671w1672w & wire_y_pipeff_2_w_lg_w_q_range1665w1666w & wire_y_pipeff_2_w_lg_w_q_range1659w1660w & wire_y_pipeff_2_w_lg_w_q_range1653w1654w & wire_y_pipeff_2_w_lg_w_q_range1647w1648w & wire_y_pipeff_2_w_lg_w_q_range1641w1642w & wire_y_pipeff_2_w_lg_w_q_range1635w1636w & wire_y_pipeff_2_w_lg_w_q_range1629w1630w & wire_y_pipeff_2_w_lg_w_q_range1623w1624w & wire_y_pipeff_2_w_lg_w_q_range1617w1618w & wire_y_pipeff_2_w_lg_w_q_range1611w1612w & wire_y_pipeff_2_w_lg_w_q_range1605w1606w & wire_y_pipeff_2_w_lg_w_q_range1599w1600w & wire_y_pipeff_2_w_lg_w_q_range1593w1594w & wire_y_pipeff_2_w_lg_w_q_range1587w1588w & wire_y_pipeff_2_w_lg_w_q_range1581w1582w & wire_y_pipeff_2_w_lg_w_q_range1575w1576w & wire_y_pipeff_2_w_lg_w_q_range1569w1570w & wire_y_pipeff_2_w_lg_w_q_range1563w1564w & wire_y_pipeff_2_w_lg_w_q_range1557w1558w & wire_y_pipeff_2_w_lg_w_q_range1551w1552w & wire_y_pipeff_2_w_lg_w_q_range1545w1546w & wire_y_pipeff_2_w_lg_w_q_range1539w1540w & wire_y_pipeff_2_w_lg_w_q_range1533w1534w & wire_y_pipeff_2_w_lg_w_q_range1527w1528w & wire_y_pipeff_2_w_lg_w_q_range1522w1523w);
	x_prenodeone_4_w <= ( wire_y_pipeff_3_w_lg_w_q_range2297w2298w & wire_y_pipeff_3_w_lg_w_q_range2297w2298w & wire_y_pipeff_3_w_lg_w_q_range2297w2298w & wire_y_pipeff_3_w_lg_w_q_range2297w2298w & wire_y_pipeff_3_w_lg_w_q_range2483w2484w & wire_y_pipeff_3_w_lg_w_q_range2477w2478w & wire_y_pipeff_3_w_lg_w_q_range2471w2472w & wire_y_pipeff_3_w_lg_w_q_range2465w2466w & wire_y_pipeff_3_w_lg_w_q_range2459w2460w & wire_y_pipeff_3_w_lg_w_q_range2453w2454w & wire_y_pipeff_3_w_lg_w_q_range2447w2448w & wire_y_pipeff_3_w_lg_w_q_range2441w2442w & wire_y_pipeff_3_w_lg_w_q_range2435w2436w & wire_y_pipeff_3_w_lg_w_q_range2429w2430w & wire_y_pipeff_3_w_lg_w_q_range2423w2424w & wire_y_pipeff_3_w_lg_w_q_range2417w2418w & wire_y_pipeff_3_w_lg_w_q_range2411w2412w & wire_y_pipeff_3_w_lg_w_q_range2405w2406w & wire_y_pipeff_3_w_lg_w_q_range2399w2400w & wire_y_pipeff_3_w_lg_w_q_range2393w2394w & wire_y_pipeff_3_w_lg_w_q_range2387w2388w & wire_y_pipeff_3_w_lg_w_q_range2381w2382w & wire_y_pipeff_3_w_lg_w_q_range2375w2376w & wire_y_pipeff_3_w_lg_w_q_range2369w2370w & wire_y_pipeff_3_w_lg_w_q_range2363w2364w & wire_y_pipeff_3_w_lg_w_q_range2357w2358w & wire_y_pipeff_3_w_lg_w_q_range2351w2352w & wire_y_pipeff_3_w_lg_w_q_range2345w2346w & wire_y_pipeff_3_w_lg_w_q_range2339w2340w & wire_y_pipeff_3_w_lg_w_q_range2333w2334w & wire_y_pipeff_3_w_lg_w_q_range2327w2328w & wire_y_pipeff_3_w_lg_w_q_range2322w2323w);
	x_prenodeone_5_w <= ( wire_y_pipeff_4_w_lg_w_q_range3088w3089w & wire_y_pipeff_4_w_lg_w_q_range3088w3089w & wire_y_pipeff_4_w_lg_w_q_range3088w3089w & wire_y_pipeff_4_w_lg_w_q_range3088w3089w & wire_y_pipeff_4_w_lg_w_q_range3088w3089w & wire_y_pipeff_4_w_lg_w_q_range3272w3273w & wire_y_pipeff_4_w_lg_w_q_range3266w3267w & wire_y_pipeff_4_w_lg_w_q_range3260w3261w & wire_y_pipeff_4_w_lg_w_q_range3254w3255w & wire_y_pipeff_4_w_lg_w_q_range3248w3249w & wire_y_pipeff_4_w_lg_w_q_range3242w3243w & wire_y_pipeff_4_w_lg_w_q_range3236w3237w & wire_y_pipeff_4_w_lg_w_q_range3230w3231w & wire_y_pipeff_4_w_lg_w_q_range3224w3225w & wire_y_pipeff_4_w_lg_w_q_range3218w3219w & wire_y_pipeff_4_w_lg_w_q_range3212w3213w & wire_y_pipeff_4_w_lg_w_q_range3206w3207w & wire_y_pipeff_4_w_lg_w_q_range3200w3201w & wire_y_pipeff_4_w_lg_w_q_range3194w3195w & wire_y_pipeff_4_w_lg_w_q_range3188w3189w & wire_y_pipeff_4_w_lg_w_q_range3182w3183w & wire_y_pipeff_4_w_lg_w_q_range3176w3177w & wire_y_pipeff_4_w_lg_w_q_range3170w3171w & wire_y_pipeff_4_w_lg_w_q_range3164w3165w & wire_y_pipeff_4_w_lg_w_q_range3158w3159w & wire_y_pipeff_4_w_lg_w_q_range3152w3153w & wire_y_pipeff_4_w_lg_w_q_range3146w3147w & wire_y_pipeff_4_w_lg_w_q_range3140w3141w & wire_y_pipeff_4_w_lg_w_q_range3134w3135w & wire_y_pipeff_4_w_lg_w_q_range3128w3129w & wire_y_pipeff_4_w_lg_w_q_range3122w3123w & wire_y_pipeff_4_w_lg_w_q_range3117w3118w);
	x_prenodeone_6_w <= ( wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range4056w4057w & wire_y_pipeff_5_w_lg_w_q_range4050w4051w & wire_y_pipeff_5_w_lg_w_q_range4044w4045w & wire_y_pipeff_5_w_lg_w_q_range4038w4039w & wire_y_pipeff_5_w_lg_w_q_range4032w4033w & wire_y_pipeff_5_w_lg_w_q_range4026w4027w & wire_y_pipeff_5_w_lg_w_q_range4020w4021w & wire_y_pipeff_5_w_lg_w_q_range4014w4015w & wire_y_pipeff_5_w_lg_w_q_range4008w4009w & wire_y_pipeff_5_w_lg_w_q_range4002w4003w & wire_y_pipeff_5_w_lg_w_q_range3996w3997w & wire_y_pipeff_5_w_lg_w_q_range3990w3991w & wire_y_pipeff_5_w_lg_w_q_range3984w3985w & wire_y_pipeff_5_w_lg_w_q_range3978w3979w & wire_y_pipeff_5_w_lg_w_q_range3972w3973w & wire_y_pipeff_5_w_lg_w_q_range3966w3967w & wire_y_pipeff_5_w_lg_w_q_range3960w3961w & wire_y_pipeff_5_w_lg_w_q_range3954w3955w & wire_y_pipeff_5_w_lg_w_q_range3948w3949w & wire_y_pipeff_5_w_lg_w_q_range3942w3943w & wire_y_pipeff_5_w_lg_w_q_range3936w3937w & wire_y_pipeff_5_w_lg_w_q_range3930w3931w & wire_y_pipeff_5_w_lg_w_q_range3924w3925w & wire_y_pipeff_5_w_lg_w_q_range3918w3919w & wire_y_pipeff_5_w_lg_w_q_range3912w3913w & wire_y_pipeff_5_w_lg_w_q_range3907w3908w);
	x_prenodeone_7_w <= ( wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4835w4836w & wire_y_pipeff_6_w_lg_w_q_range4829w4830w & wire_y_pipeff_6_w_lg_w_q_range4823w4824w & wire_y_pipeff_6_w_lg_w_q_range4817w4818w & wire_y_pipeff_6_w_lg_w_q_range4811w4812w & wire_y_pipeff_6_w_lg_w_q_range4805w4806w & wire_y_pipeff_6_w_lg_w_q_range4799w4800w & wire_y_pipeff_6_w_lg_w_q_range4793w4794w & wire_y_pipeff_6_w_lg_w_q_range4787w4788w & wire_y_pipeff_6_w_lg_w_q_range4781w4782w & wire_y_pipeff_6_w_lg_w_q_range4775w4776w & wire_y_pipeff_6_w_lg_w_q_range4769w4770w & wire_y_pipeff_6_w_lg_w_q_range4763w4764w & wire_y_pipeff_6_w_lg_w_q_range4757w4758w & wire_y_pipeff_6_w_lg_w_q_range4751w4752w & wire_y_pipeff_6_w_lg_w_q_range4745w4746w & wire_y_pipeff_6_w_lg_w_q_range4739w4740w & wire_y_pipeff_6_w_lg_w_q_range4733w4734w & wire_y_pipeff_6_w_lg_w_q_range4727w4728w & wire_y_pipeff_6_w_lg_w_q_range4721w4722w & wire_y_pipeff_6_w_lg_w_q_range4715w4716w & wire_y_pipeff_6_w_lg_w_q_range4709w4710w & wire_y_pipeff_6_w_lg_w_q_range4703w4704w & wire_y_pipeff_6_w_lg_w_q_range4697w4698w & wire_y_pipeff_6_w_lg_w_q_range4692w4693w);
	x_prenodeone_8_w <= ( wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5609w5610w & wire_y_pipeff_7_w_lg_w_q_range5603w5604w & wire_y_pipeff_7_w_lg_w_q_range5597w5598w & wire_y_pipeff_7_w_lg_w_q_range5591w5592w & wire_y_pipeff_7_w_lg_w_q_range5585w5586w & wire_y_pipeff_7_w_lg_w_q_range5579w5580w & wire_y_pipeff_7_w_lg_w_q_range5573w5574w & wire_y_pipeff_7_w_lg_w_q_range5567w5568w & wire_y_pipeff_7_w_lg_w_q_range5561w5562w & wire_y_pipeff_7_w_lg_w_q_range5555w5556w & wire_y_pipeff_7_w_lg_w_q_range5549w5550w & wire_y_pipeff_7_w_lg_w_q_range5543w5544w & wire_y_pipeff_7_w_lg_w_q_range5537w5538w & wire_y_pipeff_7_w_lg_w_q_range5531w5532w & wire_y_pipeff_7_w_lg_w_q_range5525w5526w & wire_y_pipeff_7_w_lg_w_q_range5519w5520w & wire_y_pipeff_7_w_lg_w_q_range5513w5514w & wire_y_pipeff_7_w_lg_w_q_range5507w5508w & wire_y_pipeff_7_w_lg_w_q_range5501w5502w & wire_y_pipeff_7_w_lg_w_q_range5495w5496w & wire_y_pipeff_7_w_lg_w_q_range5489w5490w & wire_y_pipeff_7_w_lg_w_q_range5483w5484w & wire_y_pipeff_7_w_lg_w_q_range5477w5478w & wire_y_pipeff_7_w_lg_w_q_range5472w5473w);
	x_prenodeone_9_w <= ( wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6378w6379w & wire_y_pipeff_8_w_lg_w_q_range6372w6373w & wire_y_pipeff_8_w_lg_w_q_range6366w6367w & wire_y_pipeff_8_w_lg_w_q_range6360w6361w & wire_y_pipeff_8_w_lg_w_q_range6354w6355w & wire_y_pipeff_8_w_lg_w_q_range6348w6349w & wire_y_pipeff_8_w_lg_w_q_range6342w6343w & wire_y_pipeff_8_w_lg_w_q_range6336w6337w & wire_y_pipeff_8_w_lg_w_q_range6330w6331w & wire_y_pipeff_8_w_lg_w_q_range6324w6325w & wire_y_pipeff_8_w_lg_w_q_range6318w6319w & wire_y_pipeff_8_w_lg_w_q_range6312w6313w & wire_y_pipeff_8_w_lg_w_q_range6306w6307w & wire_y_pipeff_8_w_lg_w_q_range6300w6301w & wire_y_pipeff_8_w_lg_w_q_range6294w6295w & wire_y_pipeff_8_w_lg_w_q_range6288w6289w & wire_y_pipeff_8_w_lg_w_q_range6282w6283w & wire_y_pipeff_8_w_lg_w_q_range6276w6277w & wire_y_pipeff_8_w_lg_w_q_range6270w6271w & wire_y_pipeff_8_w_lg_w_q_range6264w6265w & wire_y_pipeff_8_w_lg_w_q_range6258w6259w & wire_y_pipeff_8_w_lg_w_q_range6252w6253w & wire_y_pipeff_8_w_lg_w_q_range6247w6248w);
	x_prenodetwo_10_w <= ( wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range6968w6969w & wire_y_pipeff_9_w_lg_w_q_range7142w7143w & wire_y_pipeff_9_w_lg_w_q_range7136w7137w & wire_y_pipeff_9_w_lg_w_q_range7130w7131w & wire_y_pipeff_9_w_lg_w_q_range7124w7125w & wire_y_pipeff_9_w_lg_w_q_range7118w7119w & wire_y_pipeff_9_w_lg_w_q_range7112w7113w & wire_y_pipeff_9_w_lg_w_q_range7106w7107w & wire_y_pipeff_9_w_lg_w_q_range7100w7101w & wire_y_pipeff_9_w_lg_w_q_range7094w7095w & wire_y_pipeff_9_w_lg_w_q_range7088w7089w & wire_y_pipeff_9_w_lg_w_q_range7082w7083w & wire_y_pipeff_9_w_lg_w_q_range7076w7077w & wire_y_pipeff_9_w_lg_w_q_range7070w7071w & wire_y_pipeff_9_w_lg_w_q_range7064w7065w & wire_y_pipeff_9_w_lg_w_q_range7058w7059w & wire_y_pipeff_9_w_lg_w_q_range7052w7053w & wire_y_pipeff_9_w_lg_w_q_range7046w7047w & wire_y_pipeff_9_w_lg_w_q_range7040w7041w & wire_y_pipeff_9_w_lg_w_q_range7034w7035w);
	x_prenodetwo_11_w <= ( wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7729w7730w & wire_y_pipeff_10_w_lg_w_q_range7901w7902w & wire_y_pipeff_10_w_lg_w_q_range7895w7896w & wire_y_pipeff_10_w_lg_w_q_range7889w7890w & wire_y_pipeff_10_w_lg_w_q_range7883w7884w & wire_y_pipeff_10_w_lg_w_q_range7877w7878w & wire_y_pipeff_10_w_lg_w_q_range7871w7872w & wire_y_pipeff_10_w_lg_w_q_range7865w7866w & wire_y_pipeff_10_w_lg_w_q_range7859w7860w & wire_y_pipeff_10_w_lg_w_q_range7853w7854w & wire_y_pipeff_10_w_lg_w_q_range7847w7848w & wire_y_pipeff_10_w_lg_w_q_range7841w7842w & wire_y_pipeff_10_w_lg_w_q_range7835w7836w & wire_y_pipeff_10_w_lg_w_q_range7829w7830w & wire_y_pipeff_10_w_lg_w_q_range7823w7824w & wire_y_pipeff_10_w_lg_w_q_range7817w7818w & wire_y_pipeff_10_w_lg_w_q_range7811w7812w & wire_y_pipeff_10_w_lg_w_q_range7805w7806w & wire_y_pipeff_10_w_lg_w_q_range7799w7800w);
	x_prenodetwo_12_w <= ( wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8485w8486w & wire_y_pipeff_11_w_lg_w_q_range8655w8656w & wire_y_pipeff_11_w_lg_w_q_range8649w8650w & wire_y_pipeff_11_w_lg_w_q_range8643w8644w & wire_y_pipeff_11_w_lg_w_q_range8637w8638w & wire_y_pipeff_11_w_lg_w_q_range8631w8632w & wire_y_pipeff_11_w_lg_w_q_range8625w8626w & wire_y_pipeff_11_w_lg_w_q_range8619w8620w & wire_y_pipeff_11_w_lg_w_q_range8613w8614w & wire_y_pipeff_11_w_lg_w_q_range8607w8608w & wire_y_pipeff_11_w_lg_w_q_range8601w8602w & wire_y_pipeff_11_w_lg_w_q_range8595w8596w & wire_y_pipeff_11_w_lg_w_q_range8589w8590w & wire_y_pipeff_11_w_lg_w_q_range8583w8584w & wire_y_pipeff_11_w_lg_w_q_range8577w8578w & wire_y_pipeff_11_w_lg_w_q_range8571w8572w & wire_y_pipeff_11_w_lg_w_q_range8565w8566w & wire_y_pipeff_11_w_lg_w_q_range8559w8560w);
	x_prenodetwo_13_w <= ( wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9236w9237w & wire_y_pipeff_12_w_lg_w_q_range9404w9405w & wire_y_pipeff_12_w_lg_w_q_range9398w9399w & wire_y_pipeff_12_w_lg_w_q_range9392w9393w & wire_y_pipeff_12_w_lg_w_q_range9386w9387w & wire_y_pipeff_12_w_lg_w_q_range9380w9381w & wire_y_pipeff_12_w_lg_w_q_range9374w9375w & wire_y_pipeff_12_w_lg_w_q_range9368w9369w & wire_y_pipeff_12_w_lg_w_q_range9362w9363w & wire_y_pipeff_12_w_lg_w_q_range9356w9357w & wire_y_pipeff_12_w_lg_w_q_range9350w9351w & wire_y_pipeff_12_w_lg_w_q_range9344w9345w & wire_y_pipeff_12_w_lg_w_q_range9338w9339w & wire_y_pipeff_12_w_lg_w_q_range9332w9333w & wire_y_pipeff_12_w_lg_w_q_range9326w9327w & wire_y_pipeff_12_w_lg_w_q_range9320w9321w & wire_y_pipeff_12_w_lg_w_q_range9314w9315w);
	x_prenodetwo_2_w <= ( wire_y_pipeff_1_w_lg_w_q_range700w701w & wire_y_pipeff_1_w_lg_w_q_range700w701w & wire_y_pipeff_1_w_lg_w_q_range700w701w & wire_y_pipeff_1_w_lg_w_q_range700w701w & wire_y_pipeff_1_w_lg_w_q_range700w701w & wire_y_pipeff_1_w_lg_w_q_range890w891w & wire_y_pipeff_1_w_lg_w_q_range884w885w & wire_y_pipeff_1_w_lg_w_q_range878w879w & wire_y_pipeff_1_w_lg_w_q_range872w873w & wire_y_pipeff_1_w_lg_w_q_range866w867w & wire_y_pipeff_1_w_lg_w_q_range860w861w & wire_y_pipeff_1_w_lg_w_q_range854w855w & wire_y_pipeff_1_w_lg_w_q_range848w849w & wire_y_pipeff_1_w_lg_w_q_range842w843w & wire_y_pipeff_1_w_lg_w_q_range836w837w & wire_y_pipeff_1_w_lg_w_q_range830w831w & wire_y_pipeff_1_w_lg_w_q_range824w825w & wire_y_pipeff_1_w_lg_w_q_range818w819w & wire_y_pipeff_1_w_lg_w_q_range812w813w & wire_y_pipeff_1_w_lg_w_q_range806w807w & wire_y_pipeff_1_w_lg_w_q_range800w801w & wire_y_pipeff_1_w_lg_w_q_range794w795w & wire_y_pipeff_1_w_lg_w_q_range788w789w & wire_y_pipeff_1_w_lg_w_q_range782w783w & wire_y_pipeff_1_w_lg_w_q_range776w777w & wire_y_pipeff_1_w_lg_w_q_range770w771w & wire_y_pipeff_1_w_lg_w_q_range764w765w & wire_y_pipeff_1_w_lg_w_q_range758w759w & wire_y_pipeff_1_w_lg_w_q_range752w753w & wire_y_pipeff_1_w_lg_w_q_range746w747w & wire_y_pipeff_1_w_lg_w_q_range740w741w & wire_y_pipeff_1_w_lg_w_q_range734w735w);
	x_prenodetwo_3_w <= ( wire_y_pipeff_2_w_lg_w_q_range1501w1502w & wire_y_pipeff_2_w_lg_w_q_range1501w1502w & wire_y_pipeff_2_w_lg_w_q_range1501w1502w & wire_y_pipeff_2_w_lg_w_q_range1501w1502w & wire_y_pipeff_2_w_lg_w_q_range1501w1502w & wire_y_pipeff_2_w_lg_w_q_range1501w1502w & wire_y_pipeff_2_w_lg_w_q_range1689w1690w & wire_y_pipeff_2_w_lg_w_q_range1683w1684w & wire_y_pipeff_2_w_lg_w_q_range1677w1678w & wire_y_pipeff_2_w_lg_w_q_range1671w1672w & wire_y_pipeff_2_w_lg_w_q_range1665w1666w & wire_y_pipeff_2_w_lg_w_q_range1659w1660w & wire_y_pipeff_2_w_lg_w_q_range1653w1654w & wire_y_pipeff_2_w_lg_w_q_range1647w1648w & wire_y_pipeff_2_w_lg_w_q_range1641w1642w & wire_y_pipeff_2_w_lg_w_q_range1635w1636w & wire_y_pipeff_2_w_lg_w_q_range1629w1630w & wire_y_pipeff_2_w_lg_w_q_range1623w1624w & wire_y_pipeff_2_w_lg_w_q_range1617w1618w & wire_y_pipeff_2_w_lg_w_q_range1611w1612w & wire_y_pipeff_2_w_lg_w_q_range1605w1606w & wire_y_pipeff_2_w_lg_w_q_range1599w1600w & wire_y_pipeff_2_w_lg_w_q_range1593w1594w & wire_y_pipeff_2_w_lg_w_q_range1587w1588w & wire_y_pipeff_2_w_lg_w_q_range1581w1582w & wire_y_pipeff_2_w_lg_w_q_range1575w1576w & wire_y_pipeff_2_w_lg_w_q_range1569w1570w & wire_y_pipeff_2_w_lg_w_q_range1563w1564w & wire_y_pipeff_2_w_lg_w_q_range1557w1558w & wire_y_pipeff_2_w_lg_w_q_range1551w1552w & wire_y_pipeff_2_w_lg_w_q_range1545w1546w & wire_y_pipeff_2_w_lg_w_q_range1539w1540w);
	x_prenodetwo_4_w <= ( wire_y_pipeff_3_w_lg_w_q_range2297w2298w & wire_y_pipeff_3_w_lg_w_q_range2297w2298w & wire_y_pipeff_3_w_lg_w_q_range2297w2298w & wire_y_pipeff_3_w_lg_w_q_range2297w2298w & wire_y_pipeff_3_w_lg_w_q_range2297w2298w & wire_y_pipeff_3_w_lg_w_q_range2297w2298w & wire_y_pipeff_3_w_lg_w_q_range2297w2298w & wire_y_pipeff_3_w_lg_w_q_range2483w2484w & wire_y_pipeff_3_w_lg_w_q_range2477w2478w & wire_y_pipeff_3_w_lg_w_q_range2471w2472w & wire_y_pipeff_3_w_lg_w_q_range2465w2466w & wire_y_pipeff_3_w_lg_w_q_range2459w2460w & wire_y_pipeff_3_w_lg_w_q_range2453w2454w & wire_y_pipeff_3_w_lg_w_q_range2447w2448w & wire_y_pipeff_3_w_lg_w_q_range2441w2442w & wire_y_pipeff_3_w_lg_w_q_range2435w2436w & wire_y_pipeff_3_w_lg_w_q_range2429w2430w & wire_y_pipeff_3_w_lg_w_q_range2423w2424w & wire_y_pipeff_3_w_lg_w_q_range2417w2418w & wire_y_pipeff_3_w_lg_w_q_range2411w2412w & wire_y_pipeff_3_w_lg_w_q_range2405w2406w & wire_y_pipeff_3_w_lg_w_q_range2399w2400w & wire_y_pipeff_3_w_lg_w_q_range2393w2394w & wire_y_pipeff_3_w_lg_w_q_range2387w2388w & wire_y_pipeff_3_w_lg_w_q_range2381w2382w & wire_y_pipeff_3_w_lg_w_q_range2375w2376w & wire_y_pipeff_3_w_lg_w_q_range2369w2370w & wire_y_pipeff_3_w_lg_w_q_range2363w2364w & wire_y_pipeff_3_w_lg_w_q_range2357w2358w & wire_y_pipeff_3_w_lg_w_q_range2351w2352w & wire_y_pipeff_3_w_lg_w_q_range2345w2346w & wire_y_pipeff_3_w_lg_w_q_range2339w2340w);
	x_prenodetwo_5_w <= ( wire_y_pipeff_4_w_lg_w_q_range3088w3089w & wire_y_pipeff_4_w_lg_w_q_range3088w3089w & wire_y_pipeff_4_w_lg_w_q_range3088w3089w & wire_y_pipeff_4_w_lg_w_q_range3088w3089w & wire_y_pipeff_4_w_lg_w_q_range3088w3089w & wire_y_pipeff_4_w_lg_w_q_range3088w3089w & wire_y_pipeff_4_w_lg_w_q_range3088w3089w & wire_y_pipeff_4_w_lg_w_q_range3088w3089w & wire_y_pipeff_4_w_lg_w_q_range3272w3273w & wire_y_pipeff_4_w_lg_w_q_range3266w3267w & wire_y_pipeff_4_w_lg_w_q_range3260w3261w & wire_y_pipeff_4_w_lg_w_q_range3254w3255w & wire_y_pipeff_4_w_lg_w_q_range3248w3249w & wire_y_pipeff_4_w_lg_w_q_range3242w3243w & wire_y_pipeff_4_w_lg_w_q_range3236w3237w & wire_y_pipeff_4_w_lg_w_q_range3230w3231w & wire_y_pipeff_4_w_lg_w_q_range3224w3225w & wire_y_pipeff_4_w_lg_w_q_range3218w3219w & wire_y_pipeff_4_w_lg_w_q_range3212w3213w & wire_y_pipeff_4_w_lg_w_q_range3206w3207w & wire_y_pipeff_4_w_lg_w_q_range3200w3201w & wire_y_pipeff_4_w_lg_w_q_range3194w3195w & wire_y_pipeff_4_w_lg_w_q_range3188w3189w & wire_y_pipeff_4_w_lg_w_q_range3182w3183w & wire_y_pipeff_4_w_lg_w_q_range3176w3177w & wire_y_pipeff_4_w_lg_w_q_range3170w3171w & wire_y_pipeff_4_w_lg_w_q_range3164w3165w & wire_y_pipeff_4_w_lg_w_q_range3158w3159w & wire_y_pipeff_4_w_lg_w_q_range3152w3153w & wire_y_pipeff_4_w_lg_w_q_range3146w3147w & wire_y_pipeff_4_w_lg_w_q_range3140w3141w & wire_y_pipeff_4_w_lg_w_q_range3134w3135w);
	x_prenodetwo_6_w <= ( wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range3874w3875w & wire_y_pipeff_5_w_lg_w_q_range4056w4057w & wire_y_pipeff_5_w_lg_w_q_range4050w4051w & wire_y_pipeff_5_w_lg_w_q_range4044w4045w & wire_y_pipeff_5_w_lg_w_q_range4038w4039w & wire_y_pipeff_5_w_lg_w_q_range4032w4033w & wire_y_pipeff_5_w_lg_w_q_range4026w4027w & wire_y_pipeff_5_w_lg_w_q_range4020w4021w & wire_y_pipeff_5_w_lg_w_q_range4014w4015w & wire_y_pipeff_5_w_lg_w_q_range4008w4009w & wire_y_pipeff_5_w_lg_w_q_range4002w4003w & wire_y_pipeff_5_w_lg_w_q_range3996w3997w & wire_y_pipeff_5_w_lg_w_q_range3990w3991w & wire_y_pipeff_5_w_lg_w_q_range3984w3985w & wire_y_pipeff_5_w_lg_w_q_range3978w3979w & wire_y_pipeff_5_w_lg_w_q_range3972w3973w & wire_y_pipeff_5_w_lg_w_q_range3966w3967w & wire_y_pipeff_5_w_lg_w_q_range3960w3961w & wire_y_pipeff_5_w_lg_w_q_range3954w3955w & wire_y_pipeff_5_w_lg_w_q_range3948w3949w & wire_y_pipeff_5_w_lg_w_q_range3942w3943w & wire_y_pipeff_5_w_lg_w_q_range3936w3937w & wire_y_pipeff_5_w_lg_w_q_range3930w3931w & wire_y_pipeff_5_w_lg_w_q_range3924w3925w);
	x_prenodetwo_7_w <= ( wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4655w4656w & wire_y_pipeff_6_w_lg_w_q_range4835w4836w & wire_y_pipeff_6_w_lg_w_q_range4829w4830w & wire_y_pipeff_6_w_lg_w_q_range4823w4824w & wire_y_pipeff_6_w_lg_w_q_range4817w4818w & wire_y_pipeff_6_w_lg_w_q_range4811w4812w & wire_y_pipeff_6_w_lg_w_q_range4805w4806w & wire_y_pipeff_6_w_lg_w_q_range4799w4800w & wire_y_pipeff_6_w_lg_w_q_range4793w4794w & wire_y_pipeff_6_w_lg_w_q_range4787w4788w & wire_y_pipeff_6_w_lg_w_q_range4781w4782w & wire_y_pipeff_6_w_lg_w_q_range4775w4776w & wire_y_pipeff_6_w_lg_w_q_range4769w4770w & wire_y_pipeff_6_w_lg_w_q_range4763w4764w & wire_y_pipeff_6_w_lg_w_q_range4757w4758w & wire_y_pipeff_6_w_lg_w_q_range4751w4752w & wire_y_pipeff_6_w_lg_w_q_range4745w4746w & wire_y_pipeff_6_w_lg_w_q_range4739w4740w & wire_y_pipeff_6_w_lg_w_q_range4733w4734w & wire_y_pipeff_6_w_lg_w_q_range4727w4728w & wire_y_pipeff_6_w_lg_w_q_range4721w4722w & wire_y_pipeff_6_w_lg_w_q_range4715w4716w & wire_y_pipeff_6_w_lg_w_q_range4709w4710w);
	x_prenodetwo_8_w <= ( wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5431w5432w & wire_y_pipeff_7_w_lg_w_q_range5609w5610w & wire_y_pipeff_7_w_lg_w_q_range5603w5604w & wire_y_pipeff_7_w_lg_w_q_range5597w5598w & wire_y_pipeff_7_w_lg_w_q_range5591w5592w & wire_y_pipeff_7_w_lg_w_q_range5585w5586w & wire_y_pipeff_7_w_lg_w_q_range5579w5580w & wire_y_pipeff_7_w_lg_w_q_range5573w5574w & wire_y_pipeff_7_w_lg_w_q_range5567w5568w & wire_y_pipeff_7_w_lg_w_q_range5561w5562w & wire_y_pipeff_7_w_lg_w_q_range5555w5556w & wire_y_pipeff_7_w_lg_w_q_range5549w5550w & wire_y_pipeff_7_w_lg_w_q_range5543w5544w & wire_y_pipeff_7_w_lg_w_q_range5537w5538w & wire_y_pipeff_7_w_lg_w_q_range5531w5532w & wire_y_pipeff_7_w_lg_w_q_range5525w5526w & wire_y_pipeff_7_w_lg_w_q_range5519w5520w & wire_y_pipeff_7_w_lg_w_q_range5513w5514w & wire_y_pipeff_7_w_lg_w_q_range5507w5508w & wire_y_pipeff_7_w_lg_w_q_range5501w5502w & wire_y_pipeff_7_w_lg_w_q_range5495w5496w & wire_y_pipeff_7_w_lg_w_q_range5489w5490w);
	x_prenodetwo_9_w <= ( wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6202w6203w & wire_y_pipeff_8_w_lg_w_q_range6378w6379w & wire_y_pipeff_8_w_lg_w_q_range6372w6373w & wire_y_pipeff_8_w_lg_w_q_range6366w6367w & wire_y_pipeff_8_w_lg_w_q_range6360w6361w & wire_y_pipeff_8_w_lg_w_q_range6354w6355w & wire_y_pipeff_8_w_lg_w_q_range6348w6349w & wire_y_pipeff_8_w_lg_w_q_range6342w6343w & wire_y_pipeff_8_w_lg_w_q_range6336w6337w & wire_y_pipeff_8_w_lg_w_q_range6330w6331w & wire_y_pipeff_8_w_lg_w_q_range6324w6325w & wire_y_pipeff_8_w_lg_w_q_range6318w6319w & wire_y_pipeff_8_w_lg_w_q_range6312w6313w & wire_y_pipeff_8_w_lg_w_q_range6306w6307w & wire_y_pipeff_8_w_lg_w_q_range6300w6301w & wire_y_pipeff_8_w_lg_w_q_range6294w6295w & wire_y_pipeff_8_w_lg_w_q_range6288w6289w & wire_y_pipeff_8_w_lg_w_q_range6282w6283w & wire_y_pipeff_8_w_lg_w_q_range6276w6277w & wire_y_pipeff_8_w_lg_w_q_range6270w6271w & wire_y_pipeff_8_w_lg_w_q_range6264w6265w);
	x_start_node_w <= wire_cxs_value;
	x_subnode_10_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7464w7721w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7456w7713w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7448w7705w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7440w7697w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7432w7689w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7424w7681w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7416w7673w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7408w7665w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7400w7657w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7392w7649w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7384w7641w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7376w7633w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7368w7625w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7360w7617w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7352w7609w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7344w7601w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7336w7593w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7328w7585w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7320w7577w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7312w7569w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7304w7561w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7296w7553w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7288w7545w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7280w7537w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7272w7529w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7264w7521w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7256w7513w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7248w7505w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7240w7497w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7232w7489w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7224w7481w & wire_ccc_cordic_m_w_lg_w_x_prenode_10_w_range7214w7470w);
	x_subnode_11_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8220w8477w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8212w8469w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8204w8461w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8196w8453w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8188w8445w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8180w8437w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8172w8429w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8164w8421w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8156w8413w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8148w8405w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8140w8397w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8132w8389w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8124w8381w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8116w8373w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8108w8365w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8100w8357w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8092w8349w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8084w8341w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8076w8333w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8068w8325w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8060w8317w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8052w8309w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8044w8301w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8036w8293w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8028w8285w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8020w8277w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8012w8269w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range8004w8261w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range7996w8253w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range7988w8245w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range7980w8237w & wire_ccc_cordic_m_w_lg_w_x_prenode_11_w_range7970w8226w);
	x_subnode_12_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8971w9228w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8963w9220w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8955w9212w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8947w9204w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8939w9196w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8931w9188w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8923w9180w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8915w9172w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8907w9164w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8899w9156w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8891w9148w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8883w9140w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8875w9132w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8867w9124w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8859w9116w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8851w9108w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8843w9100w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8835w9092w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8827w9084w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8819w9076w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8811w9068w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8803w9060w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8795w9052w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8787w9044w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8779w9036w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8771w9028w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8763w9020w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8755w9012w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8747w9004w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8739w8996w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8731w8988w & wire_ccc_cordic_m_w_lg_w_x_prenode_12_w_range8721w8977w);
	x_subnode_13_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9717w9974w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9709w9966w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9701w9958w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9693w9950w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9685w9942w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9677w9934w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9669w9926w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9661w9918w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9653w9910w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9645w9902w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9637w9894w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9629w9886w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9621w9878w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9613w9870w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9605w9862w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9597w9854w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9589w9846w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9581w9838w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9573w9830w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9565w9822w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9557w9814w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9549w9806w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9541w9798w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9533w9790w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9525w9782w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9517w9774w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9509w9766w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9501w9758w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9493w9750w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9485w9742w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9477w9734w & wire_ccc_cordic_m_w_lg_w_x_prenode_13_w_range9467w9723w);
	x_subnode_2_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1236w1493w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1228w1485w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1220w1477w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1212w1469w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1204w1461w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1196w1453w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1188w1445w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1180w1437w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1172w1429w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1164w1421w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1156w1413w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1148w1405w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1140w1397w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1132w1389w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1124w1381w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1116w1373w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1108w1365w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1100w1357w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1092w1349w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1084w1341w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1076w1333w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1068w1325w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1060w1317w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1052w1309w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1044w1301w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1036w1293w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1028w1285w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1020w1277w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1012w1269w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range1004w1261w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range996w1253w & wire_ccc_cordic_m_w_lg_w_x_prenode_2_w_range986w1242w);
	x_subnode_3_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2032w2289w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2024w2281w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2016w2273w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2008w2265w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range2000w2257w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1992w2249w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1984w2241w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1976w2233w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1968w2225w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1960w2217w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1952w2209w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1944w2201w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1936w2193w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1928w2185w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1920w2177w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1912w2169w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1904w2161w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1896w2153w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1888w2145w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1880w2137w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1872w2129w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1864w2121w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1856w2113w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1848w2105w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1840w2097w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1832w2089w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1824w2081w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1816w2073w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1808w2065w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1800w2057w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1792w2049w & wire_ccc_cordic_m_w_lg_w_x_prenode_3_w_range1782w2038w);
	x_subnode_4_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2823w3080w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2815w3072w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2807w3064w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2799w3056w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2791w3048w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2783w3040w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2775w3032w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2767w3024w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2759w3016w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2751w3008w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2743w3000w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2735w2992w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2727w2984w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2719w2976w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2711w2968w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2703w2960w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2695w2952w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2687w2944w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2679w2936w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2671w2928w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2663w2920w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2655w2912w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2647w2904w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2639w2896w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2631w2888w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2623w2880w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2615w2872w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2607w2864w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2599w2856w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2591w2848w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2583w2840w & wire_ccc_cordic_m_w_lg_w_x_prenode_4_w_range2573w2829w);
	x_subnode_5_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3609w3866w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3601w3858w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3593w3850w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3585w3842w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3577w3834w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3569w3826w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3561w3818w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3553w3810w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3545w3802w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3537w3794w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3529w3786w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3521w3778w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3513w3770w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3505w3762w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3497w3754w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3489w3746w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3481w3738w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3473w3730w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3465w3722w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3457w3714w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3449w3706w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3441w3698w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3433w3690w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3425w3682w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3417w3674w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3409w3666w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3401w3658w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3393w3650w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3385w3642w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3377w3634w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3369w3626w & wire_ccc_cordic_m_w_lg_w_x_prenode_5_w_range3359w3615w);
	x_subnode_6_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4390w4647w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4382w4639w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4374w4631w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4366w4623w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4358w4615w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4350w4607w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4342w4599w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4334w4591w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4326w4583w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4318w4575w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4310w4567w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4302w4559w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4294w4551w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4286w4543w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4278w4535w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4270w4527w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4262w4519w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4254w4511w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4246w4503w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4238w4495w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4230w4487w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4222w4479w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4214w4471w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4206w4463w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4198w4455w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4190w4447w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4182w4439w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4174w4431w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4166w4423w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4158w4415w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4150w4407w & wire_ccc_cordic_m_w_lg_w_x_prenode_6_w_range4140w4396w);
	x_subnode_7_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5166w5423w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5158w5415w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5150w5407w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5142w5399w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5134w5391w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5126w5383w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5118w5375w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5110w5367w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5102w5359w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5094w5351w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5086w5343w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5078w5335w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5070w5327w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5062w5319w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5054w5311w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5046w5303w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5038w5295w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5030w5287w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5022w5279w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5014w5271w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range5006w5263w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4998w5255w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4990w5247w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4982w5239w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4974w5231w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4966w5223w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4958w5215w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4950w5207w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4942w5199w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4934w5191w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4926w5183w & wire_ccc_cordic_m_w_lg_w_x_prenode_7_w_range4916w5172w);
	x_subnode_8_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5937w6194w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5929w6186w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5921w6178w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5913w6170w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5905w6162w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5897w6154w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5889w6146w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5881w6138w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5873w6130w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5865w6122w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5857w6114w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5849w6106w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5841w6098w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5833w6090w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5825w6082w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5817w6074w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5809w6066w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5801w6058w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5793w6050w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5785w6042w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5777w6034w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5769w6026w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5761w6018w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5753w6010w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5745w6002w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5737w5994w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5729w5986w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5721w5978w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5713w5970w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5705w5962w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5697w5954w & wire_ccc_cordic_m_w_lg_w_x_prenode_8_w_range5687w5943w);
	x_subnode_9_w <= ( wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6703w6960w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6695w6952w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6687w6944w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6679w6936w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6671w6928w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6663w6920w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6655w6912w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6647w6904w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6639w6896w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6631w6888w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6623w6880w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6615w6872w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6607w6864w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6599w6856w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6591w6848w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6583w6840w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6575w6832w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6567w6824w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6559w6816w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6551w6808w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6543w6800w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6535w6792w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6527w6784w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6519w6776w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6511w6768w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6503w6760w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6495w6752w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6487w6744w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6479w6736w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6471w6728w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6463w6720w & wire_ccc_cordic_m_w_lg_w_x_prenode_9_w_range6453w6709w);
	y_pipenode_10_w <= wire_y_pipenode_10_add_result;
	y_pipenode_11_w <= wire_y_pipenode_11_add_result;
	y_pipenode_12_w <= wire_y_pipenode_12_add_result;
	y_pipenode_13_w <= wire_y_pipenode_13_add_result;
	y_pipenode_2_w <= wire_y_pipenode_2_add_result;
	y_pipenode_3_w <= wire_y_pipenode_3_add_result;
	y_pipenode_4_w <= wire_y_pipenode_4_add_result;
	y_pipenode_5_w <= wire_y_pipenode_5_add_result;
	y_pipenode_6_w <= wire_y_pipenode_6_add_result;
	y_pipenode_7_w <= wire_y_pipenode_7_add_result;
	y_pipenode_8_w <= wire_y_pipenode_8_add_result;
	y_pipenode_9_w <= wire_y_pipenode_9_add_result;
	y_prenode_10_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6990w7466w7467w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6988w7458w7459w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6986w7450w7451w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6984w7442w7443w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6982w7434w7435w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6980w7426w7427w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6978w7418w7419w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6976w7410w7411w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range6973w7402w7403w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7149w7394w7395w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7146w7386w7387w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7140w7378w7379w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7134w7370w7371w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7128w7362w7363w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7122w7354w7355w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7116w7346w7347w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7110w7338w7339w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7104w7330w7331w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7098w7322w7323w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7092w7314w7315w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7086w7306w7307w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7080w7298w7299w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7074w7290w7291w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7068w7282w7283w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7062w7274w7275w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7056w7266w7267w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7050w7258w7259w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7044w7250w7251w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7038w7242w7243w
 & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7032w7234w7235w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7026w7226w7227w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_10_w_range7021w7217w7218w);
	y_prenode_11_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7753w8222w8223w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7751w8214w8215w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7749w8206w8207w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7747w8198w8199w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7745w8190w8191w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7743w8182w8183w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7741w8174w8175w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7739w8166w8167w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7737w8158w8159w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7734w8150w8151w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7908w8142w8143w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7905w8134w8135w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7899w8126w8127w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7893w8118w8119w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7887w8110w8111w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7881w8102w8103w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7875w8094w8095w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7869w8086w8087w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7863w8078w8079w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7857w8070w8071w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7851w8062w8063w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7845w8054w8055w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7839w8046w8047w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7833w8038w8039w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7827w8030w8031w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7821w8022w8023w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7815w8014w8015w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7809w8006w8007w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7803w7998w7999w
 & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7797w7990w7991w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7791w7982w7983w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_11_w_range7786w7973w7974w);
	y_prenode_12_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8511w8973w8974w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8509w8965w8966w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8507w8957w8958w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8505w8949w8950w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8503w8941w8942w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8501w8933w8934w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8499w8925w8926w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8497w8917w8918w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8495w8909w8910w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8493w8901w8902w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8490w8893w8894w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8662w8885w8886w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8659w8877w8878w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8653w8869w8870w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8647w8861w8862w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8641w8853w8854w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8635w8845w8846w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8629w8837w8838w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8623w8829w8830w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8617w8821w8822w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8611w8813w8814w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8605w8805w8806w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8599w8797w8798w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8593w8789w8790w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8587w8781w8782w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8581w8773w8774w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8575w8765w8766w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8569w8757w8758w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8563w8749w8750w
 & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8557w8741w8742w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8551w8733w8734w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_12_w_range8546w8724w8725w);
	y_prenode_13_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9264w9719w9720w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9262w9711w9712w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9260w9703w9704w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9258w9695w9696w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9256w9687w9688w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9254w9679w9680w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9252w9671w9672w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9250w9663w9664w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9248w9655w9656w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9246w9647w9648w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9244w9639w9640w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9241w9631w9632w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9411w9623w9624w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9408w9615w9616w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9402w9607w9608w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9396w9599w9600w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9390w9591w9592w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9384w9583w9584w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9378w9575w9576w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9372w9567w9568w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9366w9559w9560w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9360w9551w9552w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9354w9543w9544w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9348w9535w9536w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9342w9527w9528w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9336w9519w9520w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9330w9511w9512w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9324w9503w9504w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9318w9495w9496w
 & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9312w9487w9488w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9306w9479w9480w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_13_w_range9301w9470w9471w);
	y_prenode_2_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range705w1238w1239w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range897w1230w1231w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range894w1222w1223w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range888w1214w1215w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range882w1206w1207w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range876w1198w1199w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range870w1190w1191w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range864w1182w1183w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range858w1174w1175w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range852w1166w1167w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range846w1158w1159w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range840w1150w1151w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range834w1142w1143w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range828w1134w1135w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range822w1126w1127w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range816w1118w1119w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range810w1110w1111w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range804w1102w1103w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range798w1094w1095w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range792w1086w1087w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range786w1078w1079w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range780w1070w1071w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range774w1062w1063w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range768w1054w1055w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range762w1046w1047w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range756w1038w1039w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range750w1030w1031w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range744w1022w1023w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range738w1014w1015w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range732w1006w1007w
 & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range726w998w999w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_2_w_range721w989w990w);
	y_prenode_3_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1509w2034w2035w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1506w2026w2027w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1696w2018w2019w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1693w2010w2011w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1687w2002w2003w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1681w1994w1995w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1675w1986w1987w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1669w1978w1979w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1663w1970w1971w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1657w1962w1963w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1651w1954w1955w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1645w1946w1947w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1639w1938w1939w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1633w1930w1931w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1627w1922w1923w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1621w1914w1915w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1615w1906w1907w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1609w1898w1899w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1603w1890w1891w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1597w1882w1883w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1591w1874w1875w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1585w1866w1867w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1579w1858w1859w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1573w1850w1851w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1567w1842w1843w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1561w1834w1835w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1555w1826w1827w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1549w1818w1819w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1543w1810w1811w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1537w1802w1803w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1531w1794w1795w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_3_w_range1526w1785w1786w);
	y_prenode_4_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2307w2825w2826w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2305w2817w2818w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2302w2809w2810w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2490w2801w2802w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2487w2793w2794w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2481w2785w2786w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2475w2777w2778w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2469w2769w2770w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2463w2761w2762w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2457w2753w2754w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2451w2745w2746w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2445w2737w2738w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2439w2729w2730w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2433w2721w2722w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2427w2713w2714w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2421w2705w2706w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2415w2697w2698w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2409w2689w2690w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2403w2681w2682w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2397w2673w2674w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2391w2665w2666w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2385w2657w2658w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2379w2649w2650w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2373w2641w2642w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2367w2633w2634w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2361w2625w2626w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2355w2617w2618w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2349w2609w2610w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2343w2601w2602w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2337w2593w2594w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2331w2585w2586w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_4_w_range2326w2576w2577w);
	y_prenode_5_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3100w3611w3612w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3098w3603w3604w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3096w3595w3596w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3093w3587w3588w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3279w3579w3580w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3276w3571w3572w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3270w3563w3564w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3264w3555w3556w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3258w3547w3548w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3252w3539w3540w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3246w3531w3532w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3240w3523w3524w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3234w3515w3516w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3228w3507w3508w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3222w3499w3500w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3216w3491w3492w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3210w3483w3484w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3204w3475w3476w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3198w3467w3468w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3192w3459w3460w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3186w3451w3452w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3180w3443w3444w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3174w3435w3436w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3168w3427w3428w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3162w3419w3420w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3156w3411w3412w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3150w3403w3404w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3144w3395w3396w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3138w3387w3388w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3132w3379w3380w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3126w3371w3372w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_5_w_range3121w3362w3363w);
	y_prenode_6_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3888w4392w4393w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3886w4384w4385w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3884w4376w4377w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3882w4368w4369w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3879w4360w4361w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4063w4352w4353w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4060w4344w4345w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4054w4336w4337w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4048w4328w4329w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4042w4320w4321w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4036w4312w4313w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4030w4304w4305w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4024w4296w4297w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4018w4288w4289w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4012w4280w4281w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4006w4272w4273w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range4000w4264w4265w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3994w4256w4257w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3988w4248w4249w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3982w4240w4241w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3976w4232w4233w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3970w4224w4225w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3964w4216w4217w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3958w4208w4209w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3952w4200w4201w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3946w4192w4193w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3940w4184w4185w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3934w4176w4177w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3928w4168w4169w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3922w4160w4161w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3916w4152w4153w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_6_w_range3911w4143w4144w);
	y_prenode_7_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4671w5168w5169w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4669w5160w5161w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4667w5152w5153w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4665w5144w5145w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4663w5136w5137w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4660w5128w5129w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4842w5120w5121w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4839w5112w5113w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4833w5104w5105w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4827w5096w5097w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4821w5088w5089w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4815w5080w5081w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4809w5072w5073w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4803w5064w5065w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4797w5056w5057w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4791w5048w5049w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4785w5040w5041w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4779w5032w5033w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4773w5024w5025w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4767w5016w5017w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4761w5008w5009w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4755w5000w5001w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4749w4992w4993w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4743w4984w4985w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4737w4976w4977w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4731w4968w4969w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4725w4960w4961w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4719w4952w4953w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4713w4944w4945w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4707w4936w4937w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4701w4928w4929w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_7_w_range4696w4919w4920w);
	y_prenode_8_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5449w5939w5940w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5447w5931w5932w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5445w5923w5924w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5443w5915w5916w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5441w5907w5908w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5439w5899w5900w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5436w5891w5892w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5616w5883w5884w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5613w5875w5876w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5607w5867w5868w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5601w5859w5860w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5595w5851w5852w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5589w5843w5844w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5583w5835w5836w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5577w5827w5828w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5571w5819w5820w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5565w5811w5812w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5559w5803w5804w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5553w5795w5796w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5547w5787w5788w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5541w5779w5780w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5535w5771w5772w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5529w5763w5764w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5523w5755w5756w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5517w5747w5748w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5511w5739w5740w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5505w5731w5732w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5499w5723w5724w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5493w5715w5716w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5487w5707w5708w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5481w5699w5700w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_8_w_range5476w5690w5691w);
	y_prenode_9_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6222w6705w6706w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6220w6697w6698w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6218w6689w6690w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6216w6681w6682w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6214w6673w6674w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6212w6665w6666w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6210w6657w6658w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6207w6649w6650w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6385w6641w6642w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6382w6633w6634w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6376w6625w6626w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6370w6617w6618w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6364w6609w6610w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6358w6601w6602w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6352w6593w6594w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6346w6585w6586w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6340w6577w6578w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6334w6569w6570w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6328w6561w6562w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6322w6553w6554w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6316w6545w6546w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6310w6537w6538w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6304w6529w6530w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6298w6521w6522w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6292w6513w6514w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6286w6505w6506w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6280w6497w6498w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6274w6489w6490w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6268w6481w6482w 
& wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6262w6473w6474w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6256w6465w6466w & wire_ccc_cordic_m_w_lg_w_lg_w_y_prenodeone_9_w_range6251w6456w6457w);
	y_prenodeone_10_w <= ( x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31 DOWNTO 9));
	y_prenodeone_11_w <= ( x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31 DOWNTO 10));
	y_prenodeone_12_w <= ( x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31 DOWNTO 11));
	y_prenodeone_13_w <= ( x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31 DOWNTO 12));
	y_prenodeone_2_w <= ( x_pipeff_1(31) & x_pipeff_1(31 DOWNTO 1));
	y_prenodeone_3_w <= ( x_pipeff_2(31) & x_pipeff_2(31) & x_pipeff_2(31 DOWNTO 2));
	y_prenodeone_4_w <= ( x_pipeff_3(31) & x_pipeff_3(31) & x_pipeff_3(31) & x_pipeff_3(31 DOWNTO 3));
	y_prenodeone_5_w <= ( x_pipeff_4(31) & x_pipeff_4(31) & x_pipeff_4(31) & x_pipeff_4(31) & x_pipeff_4(31 DOWNTO 4));
	y_prenodeone_6_w <= ( x_pipeff_5(31) & x_pipeff_5(31) & x_pipeff_5(31) & x_pipeff_5(31) & x_pipeff_5(31) & x_pipeff_5(31 DOWNTO 5));
	y_prenodeone_7_w <= ( x_pipeff_6(31) & x_pipeff_6(31) & x_pipeff_6(31) & x_pipeff_6(31) & x_pipeff_6(31) & x_pipeff_6(31) & x_pipeff_6(31 DOWNTO 6));
	y_prenodeone_8_w <= ( x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31 DOWNTO 7));
	y_prenodeone_9_w <= ( x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31 DOWNTO 8));
	y_prenodetwo_10_w <= ( x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31) & x_pipeff_9(31 DOWNTO 12));
	y_prenodetwo_11_w <= ( x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31) & x_pipeff_10(31 DOWNTO 13));
	y_prenodetwo_12_w <= ( x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31) & x_pipeff_11(31 DOWNTO 14));
	y_prenodetwo_13_w <= ( x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31) & x_pipeff_12(31 DOWNTO 15));
	y_prenodetwo_2_w <= ( x_pipeff_1(31) & x_pipeff_1(31) & x_pipeff_1(31) & x_pipeff_1(31) & x_pipeff_1(31 DOWNTO 4));
	y_prenodetwo_3_w <= ( x_pipeff_2(31) & x_pipeff_2(31) & x_pipeff_2(31) & x_pipeff_2(31) & x_pipeff_2(31) & x_pipeff_2(31 DOWNTO 5));
	y_prenodetwo_4_w <= ( x_pipeff_3(31) & x_pipeff_3(31) & x_pipeff_3(31) & x_pipeff_3(31) & x_pipeff_3(31) & x_pipeff_3(31) & x_pipeff_3(31 DOWNTO 6));
	y_prenodetwo_5_w <= ( x_pipeff_4(31) & x_pipeff_4(31) & x_pipeff_4(31) & x_pipeff_4(31) & x_pipeff_4(31) & x_pipeff_4(31) & x_pipeff_4(31) & x_pipeff_4(31 DOWNTO 7));
	y_prenodetwo_6_w <= ( x_pipeff_5(31) & x_pipeff_5(31) & x_pipeff_5(31) & x_pipeff_5(31) & x_pipeff_5(31) & x_pipeff_5(31) & x_pipeff_5(31) & x_pipeff_5(31) & x_pipeff_5(31 DOWNTO 8));
	y_prenodetwo_7_w <= ( x_pipeff_6(31) & x_pipeff_6(31) & x_pipeff_6(31) & x_pipeff_6(31) & x_pipeff_6(31) & x_pipeff_6(31) & x_pipeff_6(31) & x_pipeff_6(31) & x_pipeff_6(31) & x_pipeff_6(31 DOWNTO 9));
	y_prenodetwo_8_w <= ( x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31) & x_pipeff_7(31 DOWNTO 10));
	y_prenodetwo_9_w <= ( x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31) & x_pipeff_8(31 DOWNTO 11));
	y_subnode_10_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7468w7723w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7460w7715w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7452w7707w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7444w7699w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7436w7691w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7428w7683w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7420w7675w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7412w7667w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7404w7659w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7396w7651w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7388w7643w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7380w7635w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7372w7627w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7364w7619w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7356w7611w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7348w7603w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7340w7595w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7332w7587w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7324w7579w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7316w7571w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7308w7563w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7300w7555w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7292w7547w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7284w7539w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7276w7531w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7268w7523w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7260w7515w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7252w7507w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7244w7499w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7236w7491w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7228w7483w & wire_ccc_cordic_m_w_lg_w_y_prenode_10_w_range7219w7473w);
	y_subnode_11_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8224w8479w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8216w8471w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8208w8463w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8200w8455w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8192w8447w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8184w8439w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8176w8431w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8168w8423w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8160w8415w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8152w8407w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8144w8399w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8136w8391w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8128w8383w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8120w8375w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8112w8367w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8104w8359w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8096w8351w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8088w8343w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8080w8335w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8072w8327w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8064w8319w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8056w8311w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8048w8303w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8040w8295w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8032w8287w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8024w8279w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8016w8271w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8008w8263w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range8000w8255w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range7992w8247w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range7984w8239w & wire_ccc_cordic_m_w_lg_w_y_prenode_11_w_range7975w8229w);
	y_subnode_12_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8975w9230w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8967w9222w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8959w9214w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8951w9206w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8943w9198w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8935w9190w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8927w9182w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8919w9174w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8911w9166w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8903w9158w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8895w9150w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8887w9142w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8879w9134w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8871w9126w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8863w9118w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8855w9110w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8847w9102w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8839w9094w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8831w9086w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8823w9078w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8815w9070w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8807w9062w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8799w9054w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8791w9046w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8783w9038w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8775w9030w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8767w9022w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8759w9014w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8751w9006w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8743w8998w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8735w8990w & wire_ccc_cordic_m_w_lg_w_y_prenode_12_w_range8726w8980w);
	y_subnode_13_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9721w9976w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9713w9968w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9705w9960w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9697w9952w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9689w9944w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9681w9936w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9673w9928w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9665w9920w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9657w9912w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9649w9904w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9641w9896w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9633w9888w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9625w9880w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9617w9872w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9609w9864w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9601w9856w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9593w9848w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9585w9840w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9577w9832w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9569w9824w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9561w9816w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9553w9808w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9545w9800w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9537w9792w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9529w9784w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9521w9776w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9513w9768w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9505w9760w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9497w9752w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9489w9744w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9481w9736w & wire_ccc_cordic_m_w_lg_w_y_prenode_13_w_range9472w9726w);
	y_subnode_1_w <= ( wire_x_pipeff_0_w_lg_w_q_range689w698w & wire_x_pipeff_0_w_lg_w_q_range684w696w & wire_x_pipeff_0_w_lg_w_q_range679w694w & wire_x_pipeff_0_w_lg_w_lg_w_q_range674w691w692w & wire_x_pipeff_0_w_lg_w_lg_w_q_range669w686w687w & wire_x_pipeff_0_w_lg_w_lg_w_q_range664w681w682w & wire_x_pipeff_0_w_lg_w_lg_w_q_range659w676w677w & wire_x_pipeff_0_w_lg_w_lg_w_q_range654w671w672w & wire_x_pipeff_0_w_lg_w_lg_w_q_range649w666w667w & wire_x_pipeff_0_w_lg_w_lg_w_q_range644w661w662w & wire_x_pipeff_0_w_lg_w_lg_w_q_range639w656w657w & wire_x_pipeff_0_w_lg_w_lg_w_q_range634w651w652w & wire_x_pipeff_0_w_lg_w_lg_w_q_range629w646w647w & wire_x_pipeff_0_w_lg_w_lg_w_q_range624w641w642w & wire_x_pipeff_0_w_lg_w_lg_w_q_range619w636w637w & wire_x_pipeff_0_w_lg_w_lg_w_q_range614w631w632w & wire_x_pipeff_0_w_lg_w_lg_w_q_range609w626w627w & wire_x_pipeff_0_w_lg_w_lg_w_q_range604w621w622w & wire_x_pipeff_0_w_lg_w_lg_w_q_range599w616w617w & wire_x_pipeff_0_w_lg_w_lg_w_q_range594w611w612w & wire_x_pipeff_0_w_lg_w_lg_w_q_range589w606w607w & wire_x_pipeff_0_w_lg_w_lg_w_q_range584w601w602w & wire_x_pipeff_0_w_lg_w_lg_w_q_range579w596w597w & wire_x_pipeff_0_w_lg_w_lg_w_q_range574w591w592w & wire_x_pipeff_0_w_lg_w_lg_w_q_range569w586w587w & wire_x_pipeff_0_w_lg_w_lg_w_q_range564w581w582w & wire_x_pipeff_0_w_lg_w_lg_w_q_range558w576w577w & wire_x_pipeff_0_w_lg_w_lg_w_q_range552w571w572w & wire_x_pipeff_0_w_lg_w_lg_w_q_range544w566w567w & wire_x_pipeff_0_w_lg_w_lg_w_q_range560w561w562w & wire_x_pipeff_0_w_lg_w_lg_w_q_range554w555w556w & wire_x_pipeff_0_w_lg_w_lg_w_q_range547w548w549w);
	y_subnode_2_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1240w1495w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1232w1487w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1224w1479w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1216w1471w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1208w1463w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1200w1455w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1192w1447w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1184w1439w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1176w1431w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1168w1423w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1160w1415w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1152w1407w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1144w1399w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1136w1391w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1128w1383w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1120w1375w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1112w1367w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1104w1359w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1096w1351w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1088w1343w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1080w1335w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1072w1327w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1064w1319w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1056w1311w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1048w1303w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1040w1295w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1032w1287w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1024w1279w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1016w1271w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1008w1263w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range1000w1255w & wire_ccc_cordic_m_w_lg_w_y_prenode_2_w_range991w1245w);
	y_subnode_3_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2036w2291w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2028w2283w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2020w2275w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2012w2267w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range2004w2259w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1996w2251w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1988w2243w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1980w2235w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1972w2227w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1964w2219w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1956w2211w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1948w2203w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1940w2195w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1932w2187w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1924w2179w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1916w2171w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1908w2163w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1900w2155w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1892w2147w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1884w2139w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1876w2131w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1868w2123w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1860w2115w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1852w2107w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1844w2099w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1836w2091w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1828w2083w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1820w2075w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1812w2067w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1804w2059w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1796w2051w & wire_ccc_cordic_m_w_lg_w_y_prenode_3_w_range1787w2041w);
	y_subnode_4_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2827w3082w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2819w3074w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2811w3066w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2803w3058w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2795w3050w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2787w3042w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2779w3034w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2771w3026w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2763w3018w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2755w3010w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2747w3002w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2739w2994w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2731w2986w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2723w2978w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2715w2970w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2707w2962w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2699w2954w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2691w2946w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2683w2938w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2675w2930w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2667w2922w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2659w2914w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2651w2906w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2643w2898w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2635w2890w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2627w2882w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2619w2874w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2611w2866w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2603w2858w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2595w2850w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2587w2842w & wire_ccc_cordic_m_w_lg_w_y_prenode_4_w_range2578w2832w);
	y_subnode_5_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3613w3868w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3605w3860w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3597w3852w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3589w3844w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3581w3836w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3573w3828w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3565w3820w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3557w3812w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3549w3804w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3541w3796w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3533w3788w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3525w3780w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3517w3772w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3509w3764w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3501w3756w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3493w3748w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3485w3740w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3477w3732w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3469w3724w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3461w3716w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3453w3708w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3445w3700w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3437w3692w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3429w3684w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3421w3676w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3413w3668w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3405w3660w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3397w3652w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3389w3644w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3381w3636w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3373w3628w & wire_ccc_cordic_m_w_lg_w_y_prenode_5_w_range3364w3618w);
	y_subnode_6_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4394w4649w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4386w4641w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4378w4633w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4370w4625w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4362w4617w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4354w4609w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4346w4601w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4338w4593w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4330w4585w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4322w4577w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4314w4569w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4306w4561w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4298w4553w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4290w4545w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4282w4537w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4274w4529w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4266w4521w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4258w4513w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4250w4505w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4242w4497w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4234w4489w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4226w4481w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4218w4473w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4210w4465w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4202w4457w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4194w4449w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4186w4441w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4178w4433w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4170w4425w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4162w4417w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4154w4409w & wire_ccc_cordic_m_w_lg_w_y_prenode_6_w_range4145w4399w);
	y_subnode_7_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5170w5425w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5162w5417w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5154w5409w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5146w5401w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5138w5393w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5130w5385w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5122w5377w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5114w5369w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5106w5361w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5098w5353w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5090w5345w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5082w5337w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5074w5329w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5066w5321w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5058w5313w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5050w5305w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5042w5297w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5034w5289w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5026w5281w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5018w5273w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5010w5265w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range5002w5257w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4994w5249w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4986w5241w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4978w5233w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4970w5225w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4962w5217w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4954w5209w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4946w5201w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4938w5193w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4930w5185w & wire_ccc_cordic_m_w_lg_w_y_prenode_7_w_range4921w5175w);
	y_subnode_8_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5941w6196w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5933w6188w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5925w6180w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5917w6172w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5909w6164w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5901w6156w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5893w6148w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5885w6140w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5877w6132w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5869w6124w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5861w6116w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5853w6108w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5845w6100w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5837w6092w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5829w6084w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5821w6076w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5813w6068w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5805w6060w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5797w6052w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5789w6044w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5781w6036w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5773w6028w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5765w6020w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5757w6012w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5749w6004w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5741w5996w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5733w5988w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5725w5980w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5717w5972w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5709w5964w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5701w5956w & wire_ccc_cordic_m_w_lg_w_y_prenode_8_w_range5692w5946w);
	y_subnode_9_w <= ( wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6707w6962w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6699w6954w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6691w6946w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6683w6938w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6675w6930w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6667w6922w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6659w6914w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6651w6906w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6643w6898w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6635w6890w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6627w6882w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6619w6874w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6611w6866w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6603w6858w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6595w6850w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6587w6842w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6579w6834w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6571w6826w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6563w6818w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6555w6810w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6547w6802w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6539w6794w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6531w6786w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6523w6778w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6515w6770w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6507w6762w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6499w6754w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6491w6746w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6483w6738w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6475w6730w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6467w6722w & wire_ccc_cordic_m_w_lg_w_y_prenode_9_w_range6458w6712w);
	z_pipenode_10_w <= wire_z_pipenode_10_add_result;
	z_pipenode_11_w <= wire_z_pipenode_11_add_result;
	z_pipenode_12_w <= wire_z_pipenode_12_add_result;
	z_pipenode_13_w <= wire_z_pipenode_13_add_result;
	z_pipenode_2_w <= wire_z_pipenode_2_add_result;
	z_pipenode_3_w <= wire_z_pipenode_3_add_result;
	z_pipenode_4_w <= wire_z_pipenode_4_add_result;
	z_pipenode_5_w <= wire_z_pipenode_5_add_result;
	z_pipenode_6_w <= wire_z_pipenode_6_add_result;
	z_pipenode_7_w <= wire_z_pipenode_7_add_result;
	z_pipenode_8_w <= wire_z_pipenode_8_add_result;
	z_pipenode_9_w <= wire_z_pipenode_9_add_result;
	z_subnode_10_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7725w7726w7727w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7717w7718w7719w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7709w7710w7711w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7701w7702w7703w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7693w7694w7695w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7685w7686w7687w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7677w7678w7679w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7669w7670w7671w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7661w7662w7663w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7653w7654w7655w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7645w7646w7647w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7637w7638w7639w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7629w7630w7631w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7621w7622w7623w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7613w7614w7615w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7605w7606w7607w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7597w7598w7599w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7589w7590w7591w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7581w7582w7583w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7573w7574w7575w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7565w7566w7567w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7557w7558w7559w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7549w7550w7551w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7541w7542w7543w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7533w7534w7535w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7525w7526w7527w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7517w7518w7519w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7509w7510w7511w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7501w7502w7503w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7493w7494w7495w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7485w7486w7487w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_9_w_range7476w7477w7478w);
	z_subnode_11_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8481w8482w8483w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8473w8474w8475w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8465w8466w8467w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8457w8458w8459w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8449w8450w8451w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8441w8442w8443w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8433w8434w8435w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8425w8426w8427w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8417w8418w8419w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8409w8410w8411w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8401w8402w8403w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8393w8394w8395w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8385w8386w8387w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8377w8378w8379w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8369w8370w8371w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8361w8362w8363w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8353w8354w8355w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8345w8346w8347w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8337w8338w8339w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8329w8330w8331w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8321w8322w8323w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8313w8314w8315w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8305w8306w8307w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8297w8298w8299w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8289w8290w8291w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8281w8282w8283w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8273w8274w8275w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8265w8266w8267w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8257w8258w8259w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8249w8250w8251w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8241w8242w8243w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_10_w_range8232w8233w8234w);
	z_subnode_12_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9232w9233w9234w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9224w9225w9226w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9216w9217w9218w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9208w9209w9210w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9200w9201w9202w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9192w9193w9194w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9184w9185w9186w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9176w9177w9178w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9168w9169w9170w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9160w9161w9162w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9152w9153w9154w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9144w9145w9146w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9136w9137w9138w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9128w9129w9130w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9120w9121w9122w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9112w9113w9114w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9104w9105w9106w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9096w9097w9098w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9088w9089w9090w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9080w9081w9082w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9072w9073w9074w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9064w9065w9066w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9056w9057w9058w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9048w9049w9050w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9040w9041w9042w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9032w9033w9034w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9024w9025w9026w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9016w9017w9018w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9008w9009w9010w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range9000w9001w9002w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range8992w8993w8994w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_11_w_range8983w8984w8985w);
	z_subnode_13_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9978w9979w9980w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9970w9971w9972w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9962w9963w9964w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9954w9955w9956w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9946w9947w9948w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9938w9939w9940w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9930w9931w9932w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9922w9923w9924w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9914w9915w9916w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9906w9907w9908w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9898w9899w9900w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9890w9891w9892w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9882w9883w9884w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9874w9875w9876w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9866w9867w9868w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9858w9859w9860w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9850w9851w9852w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9842w9843w9844w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9834w9835w9836w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9826w9827w9828w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9818w9819w9820w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9810w9811w9812w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9802w9803w9804w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9794w9795w9796w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9786w9787w9788w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9778w9779w9780w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9770w9771w9772w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9762w9763w9764w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9754w9755w9756w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9746w9747w9748w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9738w9739w9740w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_12_w_range9729w9730w9731w);
	z_subnode_2_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1497w1498w1499w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1489w1490w1491w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1481w1482w1483w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1473w1474w1475w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1465w1466w1467w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1457w1458w1459w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1449w1450w1451w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1441w1442w1443w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1433w1434w1435w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1425w1426w1427w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1417w1418w1419w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1409w1410w1411w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1401w1402w1403w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1393w1394w1395w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1385w1386w1387w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1377w1378w1379w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1369w1370w1371w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1361w1362w1363w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1353w1354w1355w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1345w1346w1347w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1337w1338w1339w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1329w1330w1331w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1321w1322w1323w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1313w1314w1315w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1305w1306w1307w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1297w1298w1299w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1289w1290w1291w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1281w1282w1283w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1273w1274w1275w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1265w1266w1267w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1257w1258w1259w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_1_w_range1248w1249w1250w);
	z_subnode_3_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2293w2294w2295w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2285w2286w2287w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2277w2278w2279w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2269w2270w2271w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2261w2262w2263w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2253w2254w2255w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2245w2246w2247w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2237w2238w2239w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2229w2230w2231w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2221w2222w2223w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2213w2214w2215w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2205w2206w2207w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2197w2198w2199w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2189w2190w2191w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2181w2182w2183w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2173w2174w2175w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2165w2166w2167w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2157w2158w2159w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2149w2150w2151w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2141w2142w2143w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2133w2134w2135w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2125w2126w2127w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2117w2118w2119w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2109w2110w2111w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2101w2102w2103w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2093w2094w2095w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2085w2086w2087w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2077w2078w2079w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2069w2070w2071w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2061w2062w2063w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2053w2054w2055w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_2_w_range2044w2045w2046w);
	z_subnode_4_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3084w3085w3086w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3076w3077w3078w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3068w3069w3070w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3060w3061w3062w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3052w3053w3054w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3044w3045w3046w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3036w3037w3038w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3028w3029w3030w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3020w3021w3022w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3012w3013w3014w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range3004w3005w3006w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2996w2997w2998w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2988w2989w2990w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2980w2981w2982w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2972w2973w2974w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2964w2965w2966w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2956w2957w2958w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2948w2949w2950w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2940w2941w2942w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2932w2933w2934w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2924w2925w2926w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2916w2917w2918w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2908w2909w2910w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2900w2901w2902w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2892w2893w2894w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2884w2885w2886w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2876w2877w2878w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2868w2869w2870w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2860w2861w2862w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2852w2853w2854w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2844w2845w2846w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_3_w_range2835w2836w2837w);
	z_subnode_5_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3870w3871w3872w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3862w3863w3864w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3854w3855w3856w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3846w3847w3848w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3838w3839w3840w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3830w3831w3832w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3822w3823w3824w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3814w3815w3816w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3806w3807w3808w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3798w3799w3800w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3790w3791w3792w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3782w3783w3784w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3774w3775w3776w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3766w3767w3768w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3758w3759w3760w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3750w3751w3752w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3742w3743w3744w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3734w3735w3736w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3726w3727w3728w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3718w3719w3720w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3710w3711w3712w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3702w3703w3704w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3694w3695w3696w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3686w3687w3688w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3678w3679w3680w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3670w3671w3672w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3662w3663w3664w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3654w3655w3656w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3646w3647w3648w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3638w3639w3640w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3630w3631w3632w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_4_w_range3621w3622w3623w);
	z_subnode_6_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4651w4652w4653w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4643w4644w4645w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4635w4636w4637w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4627w4628w4629w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4619w4620w4621w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4611w4612w4613w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4603w4604w4605w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4595w4596w4597w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4587w4588w4589w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4579w4580w4581w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4571w4572w4573w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4563w4564w4565w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4555w4556w4557w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4547w4548w4549w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4539w4540w4541w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4531w4532w4533w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4523w4524w4525w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4515w4516w4517w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4507w4508w4509w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4499w4500w4501w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4491w4492w4493w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4483w4484w4485w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4475w4476w4477w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4467w4468w4469w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4459w4460w4461w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4451w4452w4453w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4443w4444w4445w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4435w4436w4437w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4427w4428w4429w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4419w4420w4421w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4411w4412w4413w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_5_w_range4402w4403w4404w);
	z_subnode_7_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5427w5428w5429w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5419w5420w5421w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5411w5412w5413w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5403w5404w5405w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5395w5396w5397w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5387w5388w5389w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5379w5380w5381w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5371w5372w5373w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5363w5364w5365w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5355w5356w5357w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5347w5348w5349w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5339w5340w5341w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5331w5332w5333w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5323w5324w5325w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5315w5316w5317w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5307w5308w5309w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5299w5300w5301w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5291w5292w5293w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5283w5284w5285w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5275w5276w5277w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5267w5268w5269w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5259w5260w5261w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5251w5252w5253w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5243w5244w5245w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5235w5236w5237w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5227w5228w5229w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5219w5220w5221w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5211w5212w5213w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5203w5204w5205w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5195w5196w5197w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5187w5188w5189w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_6_w_range5178w5179w5180w);
	z_subnode_8_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6198w6199w6200w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6190w6191w6192w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6182w6183w6184w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6174w6175w6176w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6166w6167w6168w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6158w6159w6160w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6150w6151w6152w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6142w6143w6144w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6134w6135w6136w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6126w6127w6128w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6118w6119w6120w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6110w6111w6112w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6102w6103w6104w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6094w6095w6096w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6086w6087w6088w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6078w6079w6080w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6070w6071w6072w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6062w6063w6064w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6054w6055w6056w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6046w6047w6048w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6038w6039w6040w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6030w6031w6032w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6022w6023w6024w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6014w6015w6016w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range6006w6007w6008w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5998w5999w6000w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5990w5991w5992w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5982w5983w5984w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5974w5975w5976w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5966w5967w5968w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5958w5959w5960w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_7_w_range5949w5950w5951w);
	z_subnode_9_w <= ( wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6964w6965w6966w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6956w6957w6958w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6948w6949w6950w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6940w6941w6942w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6932w6933w6934w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6924w6925w6926w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6916w6917w6918w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6908w6909w6910w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6900w6901w6902w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6892w6893w6894w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6884w6885w6886w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6876w6877w6878w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6868w6869w6870w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6860w6861w6862w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6852w6853w6854w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6844w6845w6846w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6836w6837w6838w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6828w6829w6830w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6820w6821w6822w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6812w6813w6814w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6804w6805w6806w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6796w6797w6798w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6788w6789w6790w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6780w6781w6782w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6772w6773w6774w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6764w6765w6766w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6756w6757w6758w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6748w6749w6750w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6740w6741w6742w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6732w6733w6734w & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6724w6725w6726w
 & wire_ccc_cordic_m_w_lg_w_lg_w_atannode_8_w_range6715w6716w6717w);
	wire_ccc_cordic_m_w_atannode_10_w_range8232w(0) <= atannode_10_w(0);
	wire_ccc_cordic_m_w_atannode_10_w_range8313w(0) <= atannode_10_w(10);
	wire_ccc_cordic_m_w_atannode_10_w_range8321w(0) <= atannode_10_w(11);
	wire_ccc_cordic_m_w_atannode_10_w_range8329w(0) <= atannode_10_w(12);
	wire_ccc_cordic_m_w_atannode_10_w_range8337w(0) <= atannode_10_w(13);
	wire_ccc_cordic_m_w_atannode_10_w_range8345w(0) <= atannode_10_w(14);
	wire_ccc_cordic_m_w_atannode_10_w_range8353w(0) <= atannode_10_w(15);
	wire_ccc_cordic_m_w_atannode_10_w_range8361w(0) <= atannode_10_w(16);
	wire_ccc_cordic_m_w_atannode_10_w_range8369w(0) <= atannode_10_w(17);
	wire_ccc_cordic_m_w_atannode_10_w_range8377w(0) <= atannode_10_w(18);
	wire_ccc_cordic_m_w_atannode_10_w_range8385w(0) <= atannode_10_w(19);
	wire_ccc_cordic_m_w_atannode_10_w_range8241w(0) <= atannode_10_w(1);
	wire_ccc_cordic_m_w_atannode_10_w_range8393w(0) <= atannode_10_w(20);
	wire_ccc_cordic_m_w_atannode_10_w_range8401w(0) <= atannode_10_w(21);
	wire_ccc_cordic_m_w_atannode_10_w_range8409w(0) <= atannode_10_w(22);
	wire_ccc_cordic_m_w_atannode_10_w_range8417w(0) <= atannode_10_w(23);
	wire_ccc_cordic_m_w_atannode_10_w_range8425w(0) <= atannode_10_w(24);
	wire_ccc_cordic_m_w_atannode_10_w_range8433w(0) <= atannode_10_w(25);
	wire_ccc_cordic_m_w_atannode_10_w_range8441w(0) <= atannode_10_w(26);
	wire_ccc_cordic_m_w_atannode_10_w_range8449w(0) <= atannode_10_w(27);
	wire_ccc_cordic_m_w_atannode_10_w_range8457w(0) <= atannode_10_w(28);
	wire_ccc_cordic_m_w_atannode_10_w_range8465w(0) <= atannode_10_w(29);
	wire_ccc_cordic_m_w_atannode_10_w_range8249w(0) <= atannode_10_w(2);
	wire_ccc_cordic_m_w_atannode_10_w_range8473w(0) <= atannode_10_w(30);
	wire_ccc_cordic_m_w_atannode_10_w_range8481w(0) <= atannode_10_w(31);
	wire_ccc_cordic_m_w_atannode_10_w_range8257w(0) <= atannode_10_w(3);
	wire_ccc_cordic_m_w_atannode_10_w_range8265w(0) <= atannode_10_w(4);
	wire_ccc_cordic_m_w_atannode_10_w_range8273w(0) <= atannode_10_w(5);
	wire_ccc_cordic_m_w_atannode_10_w_range8281w(0) <= atannode_10_w(6);
	wire_ccc_cordic_m_w_atannode_10_w_range8289w(0) <= atannode_10_w(7);
	wire_ccc_cordic_m_w_atannode_10_w_range8297w(0) <= atannode_10_w(8);
	wire_ccc_cordic_m_w_atannode_10_w_range8305w(0) <= atannode_10_w(9);
	wire_ccc_cordic_m_w_atannode_11_w_range8983w(0) <= atannode_11_w(0);
	wire_ccc_cordic_m_w_atannode_11_w_range9064w(0) <= atannode_11_w(10);
	wire_ccc_cordic_m_w_atannode_11_w_range9072w(0) <= atannode_11_w(11);
	wire_ccc_cordic_m_w_atannode_11_w_range9080w(0) <= atannode_11_w(12);
	wire_ccc_cordic_m_w_atannode_11_w_range9088w(0) <= atannode_11_w(13);
	wire_ccc_cordic_m_w_atannode_11_w_range9096w(0) <= atannode_11_w(14);
	wire_ccc_cordic_m_w_atannode_11_w_range9104w(0) <= atannode_11_w(15);
	wire_ccc_cordic_m_w_atannode_11_w_range9112w(0) <= atannode_11_w(16);
	wire_ccc_cordic_m_w_atannode_11_w_range9120w(0) <= atannode_11_w(17);
	wire_ccc_cordic_m_w_atannode_11_w_range9128w(0) <= atannode_11_w(18);
	wire_ccc_cordic_m_w_atannode_11_w_range9136w(0) <= atannode_11_w(19);
	wire_ccc_cordic_m_w_atannode_11_w_range8992w(0) <= atannode_11_w(1);
	wire_ccc_cordic_m_w_atannode_11_w_range9144w(0) <= atannode_11_w(20);
	wire_ccc_cordic_m_w_atannode_11_w_range9152w(0) <= atannode_11_w(21);
	wire_ccc_cordic_m_w_atannode_11_w_range9160w(0) <= atannode_11_w(22);
	wire_ccc_cordic_m_w_atannode_11_w_range9168w(0) <= atannode_11_w(23);
	wire_ccc_cordic_m_w_atannode_11_w_range9176w(0) <= atannode_11_w(24);
	wire_ccc_cordic_m_w_atannode_11_w_range9184w(0) <= atannode_11_w(25);
	wire_ccc_cordic_m_w_atannode_11_w_range9192w(0) <= atannode_11_w(26);
	wire_ccc_cordic_m_w_atannode_11_w_range9200w(0) <= atannode_11_w(27);
	wire_ccc_cordic_m_w_atannode_11_w_range9208w(0) <= atannode_11_w(28);
	wire_ccc_cordic_m_w_atannode_11_w_range9216w(0) <= atannode_11_w(29);
	wire_ccc_cordic_m_w_atannode_11_w_range9000w(0) <= atannode_11_w(2);
	wire_ccc_cordic_m_w_atannode_11_w_range9224w(0) <= atannode_11_w(30);
	wire_ccc_cordic_m_w_atannode_11_w_range9232w(0) <= atannode_11_w(31);
	wire_ccc_cordic_m_w_atannode_11_w_range9008w(0) <= atannode_11_w(3);
	wire_ccc_cordic_m_w_atannode_11_w_range9016w(0) <= atannode_11_w(4);
	wire_ccc_cordic_m_w_atannode_11_w_range9024w(0) <= atannode_11_w(5);
	wire_ccc_cordic_m_w_atannode_11_w_range9032w(0) <= atannode_11_w(6);
	wire_ccc_cordic_m_w_atannode_11_w_range9040w(0) <= atannode_11_w(7);
	wire_ccc_cordic_m_w_atannode_11_w_range9048w(0) <= atannode_11_w(8);
	wire_ccc_cordic_m_w_atannode_11_w_range9056w(0) <= atannode_11_w(9);
	wire_ccc_cordic_m_w_atannode_12_w_range9729w(0) <= atannode_12_w(0);
	wire_ccc_cordic_m_w_atannode_12_w_range9810w(0) <= atannode_12_w(10);
	wire_ccc_cordic_m_w_atannode_12_w_range9818w(0) <= atannode_12_w(11);
	wire_ccc_cordic_m_w_atannode_12_w_range9826w(0) <= atannode_12_w(12);
	wire_ccc_cordic_m_w_atannode_12_w_range9834w(0) <= atannode_12_w(13);
	wire_ccc_cordic_m_w_atannode_12_w_range9842w(0) <= atannode_12_w(14);
	wire_ccc_cordic_m_w_atannode_12_w_range9850w(0) <= atannode_12_w(15);
	wire_ccc_cordic_m_w_atannode_12_w_range9858w(0) <= atannode_12_w(16);
	wire_ccc_cordic_m_w_atannode_12_w_range9866w(0) <= atannode_12_w(17);
	wire_ccc_cordic_m_w_atannode_12_w_range9874w(0) <= atannode_12_w(18);
	wire_ccc_cordic_m_w_atannode_12_w_range9882w(0) <= atannode_12_w(19);
	wire_ccc_cordic_m_w_atannode_12_w_range9738w(0) <= atannode_12_w(1);
	wire_ccc_cordic_m_w_atannode_12_w_range9890w(0) <= atannode_12_w(20);
	wire_ccc_cordic_m_w_atannode_12_w_range9898w(0) <= atannode_12_w(21);
	wire_ccc_cordic_m_w_atannode_12_w_range9906w(0) <= atannode_12_w(22);
	wire_ccc_cordic_m_w_atannode_12_w_range9914w(0) <= atannode_12_w(23);
	wire_ccc_cordic_m_w_atannode_12_w_range9922w(0) <= atannode_12_w(24);
	wire_ccc_cordic_m_w_atannode_12_w_range9930w(0) <= atannode_12_w(25);
	wire_ccc_cordic_m_w_atannode_12_w_range9938w(0) <= atannode_12_w(26);
	wire_ccc_cordic_m_w_atannode_12_w_range9946w(0) <= atannode_12_w(27);
	wire_ccc_cordic_m_w_atannode_12_w_range9954w(0) <= atannode_12_w(28);
	wire_ccc_cordic_m_w_atannode_12_w_range9962w(0) <= atannode_12_w(29);
	wire_ccc_cordic_m_w_atannode_12_w_range9746w(0) <= atannode_12_w(2);
	wire_ccc_cordic_m_w_atannode_12_w_range9970w(0) <= atannode_12_w(30);
	wire_ccc_cordic_m_w_atannode_12_w_range9978w(0) <= atannode_12_w(31);
	wire_ccc_cordic_m_w_atannode_12_w_range9754w(0) <= atannode_12_w(3);
	wire_ccc_cordic_m_w_atannode_12_w_range9762w(0) <= atannode_12_w(4);
	wire_ccc_cordic_m_w_atannode_12_w_range9770w(0) <= atannode_12_w(5);
	wire_ccc_cordic_m_w_atannode_12_w_range9778w(0) <= atannode_12_w(6);
	wire_ccc_cordic_m_w_atannode_12_w_range9786w(0) <= atannode_12_w(7);
	wire_ccc_cordic_m_w_atannode_12_w_range9794w(0) <= atannode_12_w(8);
	wire_ccc_cordic_m_w_atannode_12_w_range9802w(0) <= atannode_12_w(9);
	wire_ccc_cordic_m_w_atannode_1_w_range1248w(0) <= atannode_1_w(0);
	wire_ccc_cordic_m_w_atannode_1_w_range1329w(0) <= atannode_1_w(10);
	wire_ccc_cordic_m_w_atannode_1_w_range1337w(0) <= atannode_1_w(11);
	wire_ccc_cordic_m_w_atannode_1_w_range1345w(0) <= atannode_1_w(12);
	wire_ccc_cordic_m_w_atannode_1_w_range1353w(0) <= atannode_1_w(13);
	wire_ccc_cordic_m_w_atannode_1_w_range1361w(0) <= atannode_1_w(14);
	wire_ccc_cordic_m_w_atannode_1_w_range1369w(0) <= atannode_1_w(15);
	wire_ccc_cordic_m_w_atannode_1_w_range1377w(0) <= atannode_1_w(16);
	wire_ccc_cordic_m_w_atannode_1_w_range1385w(0) <= atannode_1_w(17);
	wire_ccc_cordic_m_w_atannode_1_w_range1393w(0) <= atannode_1_w(18);
	wire_ccc_cordic_m_w_atannode_1_w_range1401w(0) <= atannode_1_w(19);
	wire_ccc_cordic_m_w_atannode_1_w_range1257w(0) <= atannode_1_w(1);
	wire_ccc_cordic_m_w_atannode_1_w_range1409w(0) <= atannode_1_w(20);
	wire_ccc_cordic_m_w_atannode_1_w_range1417w(0) <= atannode_1_w(21);
	wire_ccc_cordic_m_w_atannode_1_w_range1425w(0) <= atannode_1_w(22);
	wire_ccc_cordic_m_w_atannode_1_w_range1433w(0) <= atannode_1_w(23);
	wire_ccc_cordic_m_w_atannode_1_w_range1441w(0) <= atannode_1_w(24);
	wire_ccc_cordic_m_w_atannode_1_w_range1449w(0) <= atannode_1_w(25);
	wire_ccc_cordic_m_w_atannode_1_w_range1457w(0) <= atannode_1_w(26);
	wire_ccc_cordic_m_w_atannode_1_w_range1465w(0) <= atannode_1_w(27);
	wire_ccc_cordic_m_w_atannode_1_w_range1473w(0) <= atannode_1_w(28);
	wire_ccc_cordic_m_w_atannode_1_w_range1481w(0) <= atannode_1_w(29);
	wire_ccc_cordic_m_w_atannode_1_w_range1265w(0) <= atannode_1_w(2);
	wire_ccc_cordic_m_w_atannode_1_w_range1489w(0) <= atannode_1_w(30);
	wire_ccc_cordic_m_w_atannode_1_w_range1497w(0) <= atannode_1_w(31);
	wire_ccc_cordic_m_w_atannode_1_w_range1273w(0) <= atannode_1_w(3);
	wire_ccc_cordic_m_w_atannode_1_w_range1281w(0) <= atannode_1_w(4);
	wire_ccc_cordic_m_w_atannode_1_w_range1289w(0) <= atannode_1_w(5);
	wire_ccc_cordic_m_w_atannode_1_w_range1297w(0) <= atannode_1_w(6);
	wire_ccc_cordic_m_w_atannode_1_w_range1305w(0) <= atannode_1_w(7);
	wire_ccc_cordic_m_w_atannode_1_w_range1313w(0) <= atannode_1_w(8);
	wire_ccc_cordic_m_w_atannode_1_w_range1321w(0) <= atannode_1_w(9);
	wire_ccc_cordic_m_w_atannode_2_w_range2044w(0) <= atannode_2_w(0);
	wire_ccc_cordic_m_w_atannode_2_w_range2125w(0) <= atannode_2_w(10);
	wire_ccc_cordic_m_w_atannode_2_w_range2133w(0) <= atannode_2_w(11);
	wire_ccc_cordic_m_w_atannode_2_w_range2141w(0) <= atannode_2_w(12);
	wire_ccc_cordic_m_w_atannode_2_w_range2149w(0) <= atannode_2_w(13);
	wire_ccc_cordic_m_w_atannode_2_w_range2157w(0) <= atannode_2_w(14);
	wire_ccc_cordic_m_w_atannode_2_w_range2165w(0) <= atannode_2_w(15);
	wire_ccc_cordic_m_w_atannode_2_w_range2173w(0) <= atannode_2_w(16);
	wire_ccc_cordic_m_w_atannode_2_w_range2181w(0) <= atannode_2_w(17);
	wire_ccc_cordic_m_w_atannode_2_w_range2189w(0) <= atannode_2_w(18);
	wire_ccc_cordic_m_w_atannode_2_w_range2197w(0) <= atannode_2_w(19);
	wire_ccc_cordic_m_w_atannode_2_w_range2053w(0) <= atannode_2_w(1);
	wire_ccc_cordic_m_w_atannode_2_w_range2205w(0) <= atannode_2_w(20);
	wire_ccc_cordic_m_w_atannode_2_w_range2213w(0) <= atannode_2_w(21);
	wire_ccc_cordic_m_w_atannode_2_w_range2221w(0) <= atannode_2_w(22);
	wire_ccc_cordic_m_w_atannode_2_w_range2229w(0) <= atannode_2_w(23);
	wire_ccc_cordic_m_w_atannode_2_w_range2237w(0) <= atannode_2_w(24);
	wire_ccc_cordic_m_w_atannode_2_w_range2245w(0) <= atannode_2_w(25);
	wire_ccc_cordic_m_w_atannode_2_w_range2253w(0) <= atannode_2_w(26);
	wire_ccc_cordic_m_w_atannode_2_w_range2261w(0) <= atannode_2_w(27);
	wire_ccc_cordic_m_w_atannode_2_w_range2269w(0) <= atannode_2_w(28);
	wire_ccc_cordic_m_w_atannode_2_w_range2277w(0) <= atannode_2_w(29);
	wire_ccc_cordic_m_w_atannode_2_w_range2061w(0) <= atannode_2_w(2);
	wire_ccc_cordic_m_w_atannode_2_w_range2285w(0) <= atannode_2_w(30);
	wire_ccc_cordic_m_w_atannode_2_w_range2293w(0) <= atannode_2_w(31);
	wire_ccc_cordic_m_w_atannode_2_w_range2069w(0) <= atannode_2_w(3);
	wire_ccc_cordic_m_w_atannode_2_w_range2077w(0) <= atannode_2_w(4);
	wire_ccc_cordic_m_w_atannode_2_w_range2085w(0) <= atannode_2_w(5);
	wire_ccc_cordic_m_w_atannode_2_w_range2093w(0) <= atannode_2_w(6);
	wire_ccc_cordic_m_w_atannode_2_w_range2101w(0) <= atannode_2_w(7);
	wire_ccc_cordic_m_w_atannode_2_w_range2109w(0) <= atannode_2_w(8);
	wire_ccc_cordic_m_w_atannode_2_w_range2117w(0) <= atannode_2_w(9);
	wire_ccc_cordic_m_w_atannode_3_w_range2835w(0) <= atannode_3_w(0);
	wire_ccc_cordic_m_w_atannode_3_w_range2916w(0) <= atannode_3_w(10);
	wire_ccc_cordic_m_w_atannode_3_w_range2924w(0) <= atannode_3_w(11);
	wire_ccc_cordic_m_w_atannode_3_w_range2932w(0) <= atannode_3_w(12);
	wire_ccc_cordic_m_w_atannode_3_w_range2940w(0) <= atannode_3_w(13);
	wire_ccc_cordic_m_w_atannode_3_w_range2948w(0) <= atannode_3_w(14);
	wire_ccc_cordic_m_w_atannode_3_w_range2956w(0) <= atannode_3_w(15);
	wire_ccc_cordic_m_w_atannode_3_w_range2964w(0) <= atannode_3_w(16);
	wire_ccc_cordic_m_w_atannode_3_w_range2972w(0) <= atannode_3_w(17);
	wire_ccc_cordic_m_w_atannode_3_w_range2980w(0) <= atannode_3_w(18);
	wire_ccc_cordic_m_w_atannode_3_w_range2988w(0) <= atannode_3_w(19);
	wire_ccc_cordic_m_w_atannode_3_w_range2844w(0) <= atannode_3_w(1);
	wire_ccc_cordic_m_w_atannode_3_w_range2996w(0) <= atannode_3_w(20);
	wire_ccc_cordic_m_w_atannode_3_w_range3004w(0) <= atannode_3_w(21);
	wire_ccc_cordic_m_w_atannode_3_w_range3012w(0) <= atannode_3_w(22);
	wire_ccc_cordic_m_w_atannode_3_w_range3020w(0) <= atannode_3_w(23);
	wire_ccc_cordic_m_w_atannode_3_w_range3028w(0) <= atannode_3_w(24);
	wire_ccc_cordic_m_w_atannode_3_w_range3036w(0) <= atannode_3_w(25);
	wire_ccc_cordic_m_w_atannode_3_w_range3044w(0) <= atannode_3_w(26);
	wire_ccc_cordic_m_w_atannode_3_w_range3052w(0) <= atannode_3_w(27);
	wire_ccc_cordic_m_w_atannode_3_w_range3060w(0) <= atannode_3_w(28);
	wire_ccc_cordic_m_w_atannode_3_w_range3068w(0) <= atannode_3_w(29);
	wire_ccc_cordic_m_w_atannode_3_w_range2852w(0) <= atannode_3_w(2);
	wire_ccc_cordic_m_w_atannode_3_w_range3076w(0) <= atannode_3_w(30);
	wire_ccc_cordic_m_w_atannode_3_w_range3084w(0) <= atannode_3_w(31);
	wire_ccc_cordic_m_w_atannode_3_w_range2860w(0) <= atannode_3_w(3);
	wire_ccc_cordic_m_w_atannode_3_w_range2868w(0) <= atannode_3_w(4);
	wire_ccc_cordic_m_w_atannode_3_w_range2876w(0) <= atannode_3_w(5);
	wire_ccc_cordic_m_w_atannode_3_w_range2884w(0) <= atannode_3_w(6);
	wire_ccc_cordic_m_w_atannode_3_w_range2892w(0) <= atannode_3_w(7);
	wire_ccc_cordic_m_w_atannode_3_w_range2900w(0) <= atannode_3_w(8);
	wire_ccc_cordic_m_w_atannode_3_w_range2908w(0) <= atannode_3_w(9);
	wire_ccc_cordic_m_w_atannode_4_w_range3621w(0) <= atannode_4_w(0);
	wire_ccc_cordic_m_w_atannode_4_w_range3702w(0) <= atannode_4_w(10);
	wire_ccc_cordic_m_w_atannode_4_w_range3710w(0) <= atannode_4_w(11);
	wire_ccc_cordic_m_w_atannode_4_w_range3718w(0) <= atannode_4_w(12);
	wire_ccc_cordic_m_w_atannode_4_w_range3726w(0) <= atannode_4_w(13);
	wire_ccc_cordic_m_w_atannode_4_w_range3734w(0) <= atannode_4_w(14);
	wire_ccc_cordic_m_w_atannode_4_w_range3742w(0) <= atannode_4_w(15);
	wire_ccc_cordic_m_w_atannode_4_w_range3750w(0) <= atannode_4_w(16);
	wire_ccc_cordic_m_w_atannode_4_w_range3758w(0) <= atannode_4_w(17);
	wire_ccc_cordic_m_w_atannode_4_w_range3766w(0) <= atannode_4_w(18);
	wire_ccc_cordic_m_w_atannode_4_w_range3774w(0) <= atannode_4_w(19);
	wire_ccc_cordic_m_w_atannode_4_w_range3630w(0) <= atannode_4_w(1);
	wire_ccc_cordic_m_w_atannode_4_w_range3782w(0) <= atannode_4_w(20);
	wire_ccc_cordic_m_w_atannode_4_w_range3790w(0) <= atannode_4_w(21);
	wire_ccc_cordic_m_w_atannode_4_w_range3798w(0) <= atannode_4_w(22);
	wire_ccc_cordic_m_w_atannode_4_w_range3806w(0) <= atannode_4_w(23);
	wire_ccc_cordic_m_w_atannode_4_w_range3814w(0) <= atannode_4_w(24);
	wire_ccc_cordic_m_w_atannode_4_w_range3822w(0) <= atannode_4_w(25);
	wire_ccc_cordic_m_w_atannode_4_w_range3830w(0) <= atannode_4_w(26);
	wire_ccc_cordic_m_w_atannode_4_w_range3838w(0) <= atannode_4_w(27);
	wire_ccc_cordic_m_w_atannode_4_w_range3846w(0) <= atannode_4_w(28);
	wire_ccc_cordic_m_w_atannode_4_w_range3854w(0) <= atannode_4_w(29);
	wire_ccc_cordic_m_w_atannode_4_w_range3638w(0) <= atannode_4_w(2);
	wire_ccc_cordic_m_w_atannode_4_w_range3862w(0) <= atannode_4_w(30);
	wire_ccc_cordic_m_w_atannode_4_w_range3870w(0) <= atannode_4_w(31);
	wire_ccc_cordic_m_w_atannode_4_w_range3646w(0) <= atannode_4_w(3);
	wire_ccc_cordic_m_w_atannode_4_w_range3654w(0) <= atannode_4_w(4);
	wire_ccc_cordic_m_w_atannode_4_w_range3662w(0) <= atannode_4_w(5);
	wire_ccc_cordic_m_w_atannode_4_w_range3670w(0) <= atannode_4_w(6);
	wire_ccc_cordic_m_w_atannode_4_w_range3678w(0) <= atannode_4_w(7);
	wire_ccc_cordic_m_w_atannode_4_w_range3686w(0) <= atannode_4_w(8);
	wire_ccc_cordic_m_w_atannode_4_w_range3694w(0) <= atannode_4_w(9);
	wire_ccc_cordic_m_w_atannode_5_w_range4402w(0) <= atannode_5_w(0);
	wire_ccc_cordic_m_w_atannode_5_w_range4483w(0) <= atannode_5_w(10);
	wire_ccc_cordic_m_w_atannode_5_w_range4491w(0) <= atannode_5_w(11);
	wire_ccc_cordic_m_w_atannode_5_w_range4499w(0) <= atannode_5_w(12);
	wire_ccc_cordic_m_w_atannode_5_w_range4507w(0) <= atannode_5_w(13);
	wire_ccc_cordic_m_w_atannode_5_w_range4515w(0) <= atannode_5_w(14);
	wire_ccc_cordic_m_w_atannode_5_w_range4523w(0) <= atannode_5_w(15);
	wire_ccc_cordic_m_w_atannode_5_w_range4531w(0) <= atannode_5_w(16);
	wire_ccc_cordic_m_w_atannode_5_w_range4539w(0) <= atannode_5_w(17);
	wire_ccc_cordic_m_w_atannode_5_w_range4547w(0) <= atannode_5_w(18);
	wire_ccc_cordic_m_w_atannode_5_w_range4555w(0) <= atannode_5_w(19);
	wire_ccc_cordic_m_w_atannode_5_w_range4411w(0) <= atannode_5_w(1);
	wire_ccc_cordic_m_w_atannode_5_w_range4563w(0) <= atannode_5_w(20);
	wire_ccc_cordic_m_w_atannode_5_w_range4571w(0) <= atannode_5_w(21);
	wire_ccc_cordic_m_w_atannode_5_w_range4579w(0) <= atannode_5_w(22);
	wire_ccc_cordic_m_w_atannode_5_w_range4587w(0) <= atannode_5_w(23);
	wire_ccc_cordic_m_w_atannode_5_w_range4595w(0) <= atannode_5_w(24);
	wire_ccc_cordic_m_w_atannode_5_w_range4603w(0) <= atannode_5_w(25);
	wire_ccc_cordic_m_w_atannode_5_w_range4611w(0) <= atannode_5_w(26);
	wire_ccc_cordic_m_w_atannode_5_w_range4619w(0) <= atannode_5_w(27);
	wire_ccc_cordic_m_w_atannode_5_w_range4627w(0) <= atannode_5_w(28);
	wire_ccc_cordic_m_w_atannode_5_w_range4635w(0) <= atannode_5_w(29);
	wire_ccc_cordic_m_w_atannode_5_w_range4419w(0) <= atannode_5_w(2);
	wire_ccc_cordic_m_w_atannode_5_w_range4643w(0) <= atannode_5_w(30);
	wire_ccc_cordic_m_w_atannode_5_w_range4651w(0) <= atannode_5_w(31);
	wire_ccc_cordic_m_w_atannode_5_w_range4427w(0) <= atannode_5_w(3);
	wire_ccc_cordic_m_w_atannode_5_w_range4435w(0) <= atannode_5_w(4);
	wire_ccc_cordic_m_w_atannode_5_w_range4443w(0) <= atannode_5_w(5);
	wire_ccc_cordic_m_w_atannode_5_w_range4451w(0) <= atannode_5_w(6);
	wire_ccc_cordic_m_w_atannode_5_w_range4459w(0) <= atannode_5_w(7);
	wire_ccc_cordic_m_w_atannode_5_w_range4467w(0) <= atannode_5_w(8);
	wire_ccc_cordic_m_w_atannode_5_w_range4475w(0) <= atannode_5_w(9);
	wire_ccc_cordic_m_w_atannode_6_w_range5178w(0) <= atannode_6_w(0);
	wire_ccc_cordic_m_w_atannode_6_w_range5259w(0) <= atannode_6_w(10);
	wire_ccc_cordic_m_w_atannode_6_w_range5267w(0) <= atannode_6_w(11);
	wire_ccc_cordic_m_w_atannode_6_w_range5275w(0) <= atannode_6_w(12);
	wire_ccc_cordic_m_w_atannode_6_w_range5283w(0) <= atannode_6_w(13);
	wire_ccc_cordic_m_w_atannode_6_w_range5291w(0) <= atannode_6_w(14);
	wire_ccc_cordic_m_w_atannode_6_w_range5299w(0) <= atannode_6_w(15);
	wire_ccc_cordic_m_w_atannode_6_w_range5307w(0) <= atannode_6_w(16);
	wire_ccc_cordic_m_w_atannode_6_w_range5315w(0) <= atannode_6_w(17);
	wire_ccc_cordic_m_w_atannode_6_w_range5323w(0) <= atannode_6_w(18);
	wire_ccc_cordic_m_w_atannode_6_w_range5331w(0) <= atannode_6_w(19);
	wire_ccc_cordic_m_w_atannode_6_w_range5187w(0) <= atannode_6_w(1);
	wire_ccc_cordic_m_w_atannode_6_w_range5339w(0) <= atannode_6_w(20);
	wire_ccc_cordic_m_w_atannode_6_w_range5347w(0) <= atannode_6_w(21);
	wire_ccc_cordic_m_w_atannode_6_w_range5355w(0) <= atannode_6_w(22);
	wire_ccc_cordic_m_w_atannode_6_w_range5363w(0) <= atannode_6_w(23);
	wire_ccc_cordic_m_w_atannode_6_w_range5371w(0) <= atannode_6_w(24);
	wire_ccc_cordic_m_w_atannode_6_w_range5379w(0) <= atannode_6_w(25);
	wire_ccc_cordic_m_w_atannode_6_w_range5387w(0) <= atannode_6_w(26);
	wire_ccc_cordic_m_w_atannode_6_w_range5395w(0) <= atannode_6_w(27);
	wire_ccc_cordic_m_w_atannode_6_w_range5403w(0) <= atannode_6_w(28);
	wire_ccc_cordic_m_w_atannode_6_w_range5411w(0) <= atannode_6_w(29);
	wire_ccc_cordic_m_w_atannode_6_w_range5195w(0) <= atannode_6_w(2);
	wire_ccc_cordic_m_w_atannode_6_w_range5419w(0) <= atannode_6_w(30);
	wire_ccc_cordic_m_w_atannode_6_w_range5427w(0) <= atannode_6_w(31);
	wire_ccc_cordic_m_w_atannode_6_w_range5203w(0) <= atannode_6_w(3);
	wire_ccc_cordic_m_w_atannode_6_w_range5211w(0) <= atannode_6_w(4);
	wire_ccc_cordic_m_w_atannode_6_w_range5219w(0) <= atannode_6_w(5);
	wire_ccc_cordic_m_w_atannode_6_w_range5227w(0) <= atannode_6_w(6);
	wire_ccc_cordic_m_w_atannode_6_w_range5235w(0) <= atannode_6_w(7);
	wire_ccc_cordic_m_w_atannode_6_w_range5243w(0) <= atannode_6_w(8);
	wire_ccc_cordic_m_w_atannode_6_w_range5251w(0) <= atannode_6_w(9);
	wire_ccc_cordic_m_w_atannode_7_w_range5949w(0) <= atannode_7_w(0);
	wire_ccc_cordic_m_w_atannode_7_w_range6030w(0) <= atannode_7_w(10);
	wire_ccc_cordic_m_w_atannode_7_w_range6038w(0) <= atannode_7_w(11);
	wire_ccc_cordic_m_w_atannode_7_w_range6046w(0) <= atannode_7_w(12);
	wire_ccc_cordic_m_w_atannode_7_w_range6054w(0) <= atannode_7_w(13);
	wire_ccc_cordic_m_w_atannode_7_w_range6062w(0) <= atannode_7_w(14);
	wire_ccc_cordic_m_w_atannode_7_w_range6070w(0) <= atannode_7_w(15);
	wire_ccc_cordic_m_w_atannode_7_w_range6078w(0) <= atannode_7_w(16);
	wire_ccc_cordic_m_w_atannode_7_w_range6086w(0) <= atannode_7_w(17);
	wire_ccc_cordic_m_w_atannode_7_w_range6094w(0) <= atannode_7_w(18);
	wire_ccc_cordic_m_w_atannode_7_w_range6102w(0) <= atannode_7_w(19);
	wire_ccc_cordic_m_w_atannode_7_w_range5958w(0) <= atannode_7_w(1);
	wire_ccc_cordic_m_w_atannode_7_w_range6110w(0) <= atannode_7_w(20);
	wire_ccc_cordic_m_w_atannode_7_w_range6118w(0) <= atannode_7_w(21);
	wire_ccc_cordic_m_w_atannode_7_w_range6126w(0) <= atannode_7_w(22);
	wire_ccc_cordic_m_w_atannode_7_w_range6134w(0) <= atannode_7_w(23);
	wire_ccc_cordic_m_w_atannode_7_w_range6142w(0) <= atannode_7_w(24);
	wire_ccc_cordic_m_w_atannode_7_w_range6150w(0) <= atannode_7_w(25);
	wire_ccc_cordic_m_w_atannode_7_w_range6158w(0) <= atannode_7_w(26);
	wire_ccc_cordic_m_w_atannode_7_w_range6166w(0) <= atannode_7_w(27);
	wire_ccc_cordic_m_w_atannode_7_w_range6174w(0) <= atannode_7_w(28);
	wire_ccc_cordic_m_w_atannode_7_w_range6182w(0) <= atannode_7_w(29);
	wire_ccc_cordic_m_w_atannode_7_w_range5966w(0) <= atannode_7_w(2);
	wire_ccc_cordic_m_w_atannode_7_w_range6190w(0) <= atannode_7_w(30);
	wire_ccc_cordic_m_w_atannode_7_w_range6198w(0) <= atannode_7_w(31);
	wire_ccc_cordic_m_w_atannode_7_w_range5974w(0) <= atannode_7_w(3);
	wire_ccc_cordic_m_w_atannode_7_w_range5982w(0) <= atannode_7_w(4);
	wire_ccc_cordic_m_w_atannode_7_w_range5990w(0) <= atannode_7_w(5);
	wire_ccc_cordic_m_w_atannode_7_w_range5998w(0) <= atannode_7_w(6);
	wire_ccc_cordic_m_w_atannode_7_w_range6006w(0) <= atannode_7_w(7);
	wire_ccc_cordic_m_w_atannode_7_w_range6014w(0) <= atannode_7_w(8);
	wire_ccc_cordic_m_w_atannode_7_w_range6022w(0) <= atannode_7_w(9);
	wire_ccc_cordic_m_w_atannode_8_w_range6715w(0) <= atannode_8_w(0);
	wire_ccc_cordic_m_w_atannode_8_w_range6796w(0) <= atannode_8_w(10);
	wire_ccc_cordic_m_w_atannode_8_w_range6804w(0) <= atannode_8_w(11);
	wire_ccc_cordic_m_w_atannode_8_w_range6812w(0) <= atannode_8_w(12);
	wire_ccc_cordic_m_w_atannode_8_w_range6820w(0) <= atannode_8_w(13);
	wire_ccc_cordic_m_w_atannode_8_w_range6828w(0) <= atannode_8_w(14);
	wire_ccc_cordic_m_w_atannode_8_w_range6836w(0) <= atannode_8_w(15);
	wire_ccc_cordic_m_w_atannode_8_w_range6844w(0) <= atannode_8_w(16);
	wire_ccc_cordic_m_w_atannode_8_w_range6852w(0) <= atannode_8_w(17);
	wire_ccc_cordic_m_w_atannode_8_w_range6860w(0) <= atannode_8_w(18);
	wire_ccc_cordic_m_w_atannode_8_w_range6868w(0) <= atannode_8_w(19);
	wire_ccc_cordic_m_w_atannode_8_w_range6724w(0) <= atannode_8_w(1);
	wire_ccc_cordic_m_w_atannode_8_w_range6876w(0) <= atannode_8_w(20);
	wire_ccc_cordic_m_w_atannode_8_w_range6884w(0) <= atannode_8_w(21);
	wire_ccc_cordic_m_w_atannode_8_w_range6892w(0) <= atannode_8_w(22);
	wire_ccc_cordic_m_w_atannode_8_w_range6900w(0) <= atannode_8_w(23);
	wire_ccc_cordic_m_w_atannode_8_w_range6908w(0) <= atannode_8_w(24);
	wire_ccc_cordic_m_w_atannode_8_w_range6916w(0) <= atannode_8_w(25);
	wire_ccc_cordic_m_w_atannode_8_w_range6924w(0) <= atannode_8_w(26);
	wire_ccc_cordic_m_w_atannode_8_w_range6932w(0) <= atannode_8_w(27);
	wire_ccc_cordic_m_w_atannode_8_w_range6940w(0) <= atannode_8_w(28);
	wire_ccc_cordic_m_w_atannode_8_w_range6948w(0) <= atannode_8_w(29);
	wire_ccc_cordic_m_w_atannode_8_w_range6732w(0) <= atannode_8_w(2);
	wire_ccc_cordic_m_w_atannode_8_w_range6956w(0) <= atannode_8_w(30);
	wire_ccc_cordic_m_w_atannode_8_w_range6964w(0) <= atannode_8_w(31);
	wire_ccc_cordic_m_w_atannode_8_w_range6740w(0) <= atannode_8_w(3);
	wire_ccc_cordic_m_w_atannode_8_w_range6748w(0) <= atannode_8_w(4);
	wire_ccc_cordic_m_w_atannode_8_w_range6756w(0) <= atannode_8_w(5);
	wire_ccc_cordic_m_w_atannode_8_w_range6764w(0) <= atannode_8_w(6);
	wire_ccc_cordic_m_w_atannode_8_w_range6772w(0) <= atannode_8_w(7);
	wire_ccc_cordic_m_w_atannode_8_w_range6780w(0) <= atannode_8_w(8);
	wire_ccc_cordic_m_w_atannode_8_w_range6788w(0) <= atannode_8_w(9);
	wire_ccc_cordic_m_w_atannode_9_w_range7476w(0) <= atannode_9_w(0);
	wire_ccc_cordic_m_w_atannode_9_w_range7557w(0) <= atannode_9_w(10);
	wire_ccc_cordic_m_w_atannode_9_w_range7565w(0) <= atannode_9_w(11);
	wire_ccc_cordic_m_w_atannode_9_w_range7573w(0) <= atannode_9_w(12);
	wire_ccc_cordic_m_w_atannode_9_w_range7581w(0) <= atannode_9_w(13);
	wire_ccc_cordic_m_w_atannode_9_w_range7589w(0) <= atannode_9_w(14);
	wire_ccc_cordic_m_w_atannode_9_w_range7597w(0) <= atannode_9_w(15);
	wire_ccc_cordic_m_w_atannode_9_w_range7605w(0) <= atannode_9_w(16);
	wire_ccc_cordic_m_w_atannode_9_w_range7613w(0) <= atannode_9_w(17);
	wire_ccc_cordic_m_w_atannode_9_w_range7621w(0) <= atannode_9_w(18);
	wire_ccc_cordic_m_w_atannode_9_w_range7629w(0) <= atannode_9_w(19);
	wire_ccc_cordic_m_w_atannode_9_w_range7485w(0) <= atannode_9_w(1);
	wire_ccc_cordic_m_w_atannode_9_w_range7637w(0) <= atannode_9_w(20);
	wire_ccc_cordic_m_w_atannode_9_w_range7645w(0) <= atannode_9_w(21);
	wire_ccc_cordic_m_w_atannode_9_w_range7653w(0) <= atannode_9_w(22);
	wire_ccc_cordic_m_w_atannode_9_w_range7661w(0) <= atannode_9_w(23);
	wire_ccc_cordic_m_w_atannode_9_w_range7669w(0) <= atannode_9_w(24);
	wire_ccc_cordic_m_w_atannode_9_w_range7677w(0) <= atannode_9_w(25);
	wire_ccc_cordic_m_w_atannode_9_w_range7685w(0) <= atannode_9_w(26);
	wire_ccc_cordic_m_w_atannode_9_w_range7693w(0) <= atannode_9_w(27);
	wire_ccc_cordic_m_w_atannode_9_w_range7701w(0) <= atannode_9_w(28);
	wire_ccc_cordic_m_w_atannode_9_w_range7709w(0) <= atannode_9_w(29);
	wire_ccc_cordic_m_w_atannode_9_w_range7493w(0) <= atannode_9_w(2);
	wire_ccc_cordic_m_w_atannode_9_w_range7717w(0) <= atannode_9_w(30);
	wire_ccc_cordic_m_w_atannode_9_w_range7725w(0) <= atannode_9_w(31);
	wire_ccc_cordic_m_w_atannode_9_w_range7501w(0) <= atannode_9_w(3);
	wire_ccc_cordic_m_w_atannode_9_w_range7509w(0) <= atannode_9_w(4);
	wire_ccc_cordic_m_w_atannode_9_w_range7517w(0) <= atannode_9_w(5);
	wire_ccc_cordic_m_w_atannode_9_w_range7525w(0) <= atannode_9_w(6);
	wire_ccc_cordic_m_w_atannode_9_w_range7533w(0) <= atannode_9_w(7);
	wire_ccc_cordic_m_w_atannode_9_w_range7541w(0) <= atannode_9_w(8);
	wire_ccc_cordic_m_w_atannode_9_w_range7549w(0) <= atannode_9_w(9);
	wire_ccc_cordic_m_w_pre_estimate_w_range9996w(0) <= pre_estimate_w(0);
	wire_ccc_cordic_m_w_pre_estimate_w_range10033w(0) <= pre_estimate_w(10);
	wire_ccc_cordic_m_w_pre_estimate_w_range10038w(0) <= pre_estimate_w(11);
	wire_ccc_cordic_m_w_pre_estimate_w_range10043w(0) <= pre_estimate_w(12);
	wire_ccc_cordic_m_w_pre_estimate_w_range10048w(0) <= pre_estimate_w(13);
	wire_ccc_cordic_m_w_pre_estimate_w_range10053w(0) <= pre_estimate_w(14);
	wire_ccc_cordic_m_w_pre_estimate_w_range10058w(0) <= pre_estimate_w(15);
	wire_ccc_cordic_m_w_pre_estimate_w_range10063w(0) <= pre_estimate_w(16);
	wire_ccc_cordic_m_w_pre_estimate_w_range10068w(0) <= pre_estimate_w(17);
	wire_ccc_cordic_m_w_pre_estimate_w_range10073w(0) <= pre_estimate_w(18);
	wire_ccc_cordic_m_w_pre_estimate_w_range10078w(0) <= pre_estimate_w(19);
	wire_ccc_cordic_m_w_pre_estimate_w_range10003w(0) <= pre_estimate_w(1);
	wire_ccc_cordic_m_w_pre_estimate_w_range10083w(0) <= pre_estimate_w(20);
	wire_ccc_cordic_m_w_pre_estimate_w_range10088w(0) <= pre_estimate_w(21);
	wire_ccc_cordic_m_w_pre_estimate_w_range10093w(0) <= pre_estimate_w(22);
	wire_ccc_cordic_m_w_pre_estimate_w_range10098w(0) <= pre_estimate_w(23);
	wire_ccc_cordic_m_w_pre_estimate_w_range10103w(0) <= pre_estimate_w(24);
	wire_ccc_cordic_m_w_pre_estimate_w_range10108w(0) <= pre_estimate_w(25);
	wire_ccc_cordic_m_w_pre_estimate_w_range10113w(0) <= pre_estimate_w(26);
	wire_ccc_cordic_m_w_pre_estimate_w_range10118w(0) <= pre_estimate_w(27);
	wire_ccc_cordic_m_w_pre_estimate_w_range10123w(0) <= pre_estimate_w(28);
	wire_ccc_cordic_m_w_pre_estimate_w_range10128w(0) <= pre_estimate_w(29);
	wire_ccc_cordic_m_w_pre_estimate_w_range10009w(0) <= pre_estimate_w(2);
	wire_ccc_cordic_m_w_pre_estimate_w_range10133w(0) <= pre_estimate_w(30);
	wire_ccc_cordic_m_w_pre_estimate_w_range10138w(0) <= pre_estimate_w(31);
	wire_ccc_cordic_m_w_pre_estimate_w_range9993w(0) <= pre_estimate_w(3);
	wire_ccc_cordic_m_w_pre_estimate_w_range10001w(0) <= pre_estimate_w(4);
	wire_ccc_cordic_m_w_pre_estimate_w_range10007w(0) <= pre_estimate_w(5);
	wire_ccc_cordic_m_w_pre_estimate_w_range10013w(0) <= pre_estimate_w(6);
	wire_ccc_cordic_m_w_pre_estimate_w_range10018w(0) <= pre_estimate_w(7);
	wire_ccc_cordic_m_w_pre_estimate_w_range10023w(0) <= pre_estimate_w(8);
	wire_ccc_cordic_m_w_pre_estimate_w_range10028w(0) <= pre_estimate_w(9);
	wire_ccc_cordic_m_w_radians_range289w(0) <= radians(0);
	wire_ccc_cordic_m_w_radians_range335w(0) <= radians(10);
	wire_ccc_cordic_m_w_radians_range340w(0) <= radians(11);
	wire_ccc_cordic_m_w_radians_range345w(0) <= radians(12);
	wire_ccc_cordic_m_w_radians_range350w(0) <= radians(13);
	wire_ccc_cordic_m_w_radians_range355w(0) <= radians(14);
	wire_ccc_cordic_m_w_radians_range360w(0) <= radians(15);
	wire_ccc_cordic_m_w_radians_range365w(0) <= radians(16);
	wire_ccc_cordic_m_w_radians_range370w(0) <= radians(17);
	wire_ccc_cordic_m_w_radians_range375w(0) <= radians(18);
	wire_ccc_cordic_m_w_radians_range380w(0) <= radians(19);
	wire_ccc_cordic_m_w_radians_range294w(0) <= radians(1);
	wire_ccc_cordic_m_w_radians_range385w(0) <= radians(20);
	wire_ccc_cordic_m_w_radians_range390w(0) <= radians(21);
	wire_ccc_cordic_m_w_radians_range395w(0) <= radians(22);
	wire_ccc_cordic_m_w_radians_range400w(0) <= radians(23);
	wire_ccc_cordic_m_w_radians_range405w(0) <= radians(24);
	wire_ccc_cordic_m_w_radians_range410w(0) <= radians(25);
	wire_ccc_cordic_m_w_radians_range415w(0) <= radians(26);
	wire_ccc_cordic_m_w_radians_range420w(0) <= radians(27);
	wire_ccc_cordic_m_w_radians_range425w(0) <= radians(28);
	wire_ccc_cordic_m_w_radians_range430w(0) <= radians(29);
	wire_ccc_cordic_m_w_radians_range297w(0) <= radians(2);
	wire_ccc_cordic_m_w_radians_range435w(0) <= radians(30);
	wire_ccc_cordic_m_w_radians_range440w(0) <= radians(31);
	wire_ccc_cordic_m_w_radians_range300w(0) <= radians(3);
	wire_ccc_cordic_m_w_radians_range305w(0) <= radians(4);
	wire_ccc_cordic_m_w_radians_range310w(0) <= radians(5);
	wire_ccc_cordic_m_w_radians_range315w(0) <= radians(6);
	wire_ccc_cordic_m_w_radians_range320w(0) <= radians(7);
	wire_ccc_cordic_m_w_radians_range325w(0) <= radians(8);
	wire_ccc_cordic_m_w_radians_range330w(0) <= radians(9);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7214w(0) <= x_prenode_10_w(0);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7296w(0) <= x_prenode_10_w(10);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7304w(0) <= x_prenode_10_w(11);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7312w(0) <= x_prenode_10_w(12);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7320w(0) <= x_prenode_10_w(13);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7328w(0) <= x_prenode_10_w(14);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7336w(0) <= x_prenode_10_w(15);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7344w(0) <= x_prenode_10_w(16);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7352w(0) <= x_prenode_10_w(17);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7360w(0) <= x_prenode_10_w(18);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7368w(0) <= x_prenode_10_w(19);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7224w(0) <= x_prenode_10_w(1);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7376w(0) <= x_prenode_10_w(20);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7384w(0) <= x_prenode_10_w(21);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7392w(0) <= x_prenode_10_w(22);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7400w(0) <= x_prenode_10_w(23);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7408w(0) <= x_prenode_10_w(24);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7416w(0) <= x_prenode_10_w(25);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7424w(0) <= x_prenode_10_w(26);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7432w(0) <= x_prenode_10_w(27);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7440w(0) <= x_prenode_10_w(28);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7448w(0) <= x_prenode_10_w(29);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7232w(0) <= x_prenode_10_w(2);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7456w(0) <= x_prenode_10_w(30);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7464w(0) <= x_prenode_10_w(31);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7240w(0) <= x_prenode_10_w(3);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7248w(0) <= x_prenode_10_w(4);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7256w(0) <= x_prenode_10_w(5);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7264w(0) <= x_prenode_10_w(6);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7272w(0) <= x_prenode_10_w(7);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7280w(0) <= x_prenode_10_w(8);
	wire_ccc_cordic_m_w_x_prenode_10_w_range7288w(0) <= x_prenode_10_w(9);
	wire_ccc_cordic_m_w_x_prenode_11_w_range7970w(0) <= x_prenode_11_w(0);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8052w(0) <= x_prenode_11_w(10);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8060w(0) <= x_prenode_11_w(11);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8068w(0) <= x_prenode_11_w(12);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8076w(0) <= x_prenode_11_w(13);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8084w(0) <= x_prenode_11_w(14);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8092w(0) <= x_prenode_11_w(15);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8100w(0) <= x_prenode_11_w(16);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8108w(0) <= x_prenode_11_w(17);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8116w(0) <= x_prenode_11_w(18);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8124w(0) <= x_prenode_11_w(19);
	wire_ccc_cordic_m_w_x_prenode_11_w_range7980w(0) <= x_prenode_11_w(1);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8132w(0) <= x_prenode_11_w(20);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8140w(0) <= x_prenode_11_w(21);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8148w(0) <= x_prenode_11_w(22);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8156w(0) <= x_prenode_11_w(23);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8164w(0) <= x_prenode_11_w(24);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8172w(0) <= x_prenode_11_w(25);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8180w(0) <= x_prenode_11_w(26);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8188w(0) <= x_prenode_11_w(27);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8196w(0) <= x_prenode_11_w(28);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8204w(0) <= x_prenode_11_w(29);
	wire_ccc_cordic_m_w_x_prenode_11_w_range7988w(0) <= x_prenode_11_w(2);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8212w(0) <= x_prenode_11_w(30);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8220w(0) <= x_prenode_11_w(31);
	wire_ccc_cordic_m_w_x_prenode_11_w_range7996w(0) <= x_prenode_11_w(3);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8004w(0) <= x_prenode_11_w(4);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8012w(0) <= x_prenode_11_w(5);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8020w(0) <= x_prenode_11_w(6);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8028w(0) <= x_prenode_11_w(7);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8036w(0) <= x_prenode_11_w(8);
	wire_ccc_cordic_m_w_x_prenode_11_w_range8044w(0) <= x_prenode_11_w(9);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8721w(0) <= x_prenode_12_w(0);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8803w(0) <= x_prenode_12_w(10);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8811w(0) <= x_prenode_12_w(11);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8819w(0) <= x_prenode_12_w(12);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8827w(0) <= x_prenode_12_w(13);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8835w(0) <= x_prenode_12_w(14);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8843w(0) <= x_prenode_12_w(15);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8851w(0) <= x_prenode_12_w(16);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8859w(0) <= x_prenode_12_w(17);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8867w(0) <= x_prenode_12_w(18);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8875w(0) <= x_prenode_12_w(19);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8731w(0) <= x_prenode_12_w(1);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8883w(0) <= x_prenode_12_w(20);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8891w(0) <= x_prenode_12_w(21);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8899w(0) <= x_prenode_12_w(22);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8907w(0) <= x_prenode_12_w(23);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8915w(0) <= x_prenode_12_w(24);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8923w(0) <= x_prenode_12_w(25);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8931w(0) <= x_prenode_12_w(26);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8939w(0) <= x_prenode_12_w(27);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8947w(0) <= x_prenode_12_w(28);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8955w(0) <= x_prenode_12_w(29);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8739w(0) <= x_prenode_12_w(2);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8963w(0) <= x_prenode_12_w(30);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8971w(0) <= x_prenode_12_w(31);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8747w(0) <= x_prenode_12_w(3);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8755w(0) <= x_prenode_12_w(4);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8763w(0) <= x_prenode_12_w(5);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8771w(0) <= x_prenode_12_w(6);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8779w(0) <= x_prenode_12_w(7);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8787w(0) <= x_prenode_12_w(8);
	wire_ccc_cordic_m_w_x_prenode_12_w_range8795w(0) <= x_prenode_12_w(9);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9467w(0) <= x_prenode_13_w(0);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9549w(0) <= x_prenode_13_w(10);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9557w(0) <= x_prenode_13_w(11);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9565w(0) <= x_prenode_13_w(12);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9573w(0) <= x_prenode_13_w(13);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9581w(0) <= x_prenode_13_w(14);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9589w(0) <= x_prenode_13_w(15);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9597w(0) <= x_prenode_13_w(16);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9605w(0) <= x_prenode_13_w(17);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9613w(0) <= x_prenode_13_w(18);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9621w(0) <= x_prenode_13_w(19);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9477w(0) <= x_prenode_13_w(1);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9629w(0) <= x_prenode_13_w(20);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9637w(0) <= x_prenode_13_w(21);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9645w(0) <= x_prenode_13_w(22);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9653w(0) <= x_prenode_13_w(23);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9661w(0) <= x_prenode_13_w(24);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9669w(0) <= x_prenode_13_w(25);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9677w(0) <= x_prenode_13_w(26);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9685w(0) <= x_prenode_13_w(27);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9693w(0) <= x_prenode_13_w(28);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9701w(0) <= x_prenode_13_w(29);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9485w(0) <= x_prenode_13_w(2);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9709w(0) <= x_prenode_13_w(30);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9717w(0) <= x_prenode_13_w(31);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9493w(0) <= x_prenode_13_w(3);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9501w(0) <= x_prenode_13_w(4);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9509w(0) <= x_prenode_13_w(5);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9517w(0) <= x_prenode_13_w(6);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9525w(0) <= x_prenode_13_w(7);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9533w(0) <= x_prenode_13_w(8);
	wire_ccc_cordic_m_w_x_prenode_13_w_range9541w(0) <= x_prenode_13_w(9);
	wire_ccc_cordic_m_w_x_prenode_2_w_range986w(0) <= x_prenode_2_w(0);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1068w(0) <= x_prenode_2_w(10);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1076w(0) <= x_prenode_2_w(11);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1084w(0) <= x_prenode_2_w(12);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1092w(0) <= x_prenode_2_w(13);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1100w(0) <= x_prenode_2_w(14);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1108w(0) <= x_prenode_2_w(15);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1116w(0) <= x_prenode_2_w(16);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1124w(0) <= x_prenode_2_w(17);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1132w(0) <= x_prenode_2_w(18);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1140w(0) <= x_prenode_2_w(19);
	wire_ccc_cordic_m_w_x_prenode_2_w_range996w(0) <= x_prenode_2_w(1);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1148w(0) <= x_prenode_2_w(20);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1156w(0) <= x_prenode_2_w(21);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1164w(0) <= x_prenode_2_w(22);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1172w(0) <= x_prenode_2_w(23);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1180w(0) <= x_prenode_2_w(24);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1188w(0) <= x_prenode_2_w(25);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1196w(0) <= x_prenode_2_w(26);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1204w(0) <= x_prenode_2_w(27);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1212w(0) <= x_prenode_2_w(28);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1220w(0) <= x_prenode_2_w(29);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1004w(0) <= x_prenode_2_w(2);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1228w(0) <= x_prenode_2_w(30);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1236w(0) <= x_prenode_2_w(31);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1012w(0) <= x_prenode_2_w(3);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1020w(0) <= x_prenode_2_w(4);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1028w(0) <= x_prenode_2_w(5);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1036w(0) <= x_prenode_2_w(6);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1044w(0) <= x_prenode_2_w(7);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1052w(0) <= x_prenode_2_w(8);
	wire_ccc_cordic_m_w_x_prenode_2_w_range1060w(0) <= x_prenode_2_w(9);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1782w(0) <= x_prenode_3_w(0);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1864w(0) <= x_prenode_3_w(10);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1872w(0) <= x_prenode_3_w(11);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1880w(0) <= x_prenode_3_w(12);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1888w(0) <= x_prenode_3_w(13);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1896w(0) <= x_prenode_3_w(14);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1904w(0) <= x_prenode_3_w(15);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1912w(0) <= x_prenode_3_w(16);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1920w(0) <= x_prenode_3_w(17);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1928w(0) <= x_prenode_3_w(18);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1936w(0) <= x_prenode_3_w(19);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1792w(0) <= x_prenode_3_w(1);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1944w(0) <= x_prenode_3_w(20);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1952w(0) <= x_prenode_3_w(21);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1960w(0) <= x_prenode_3_w(22);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1968w(0) <= x_prenode_3_w(23);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1976w(0) <= x_prenode_3_w(24);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1984w(0) <= x_prenode_3_w(25);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1992w(0) <= x_prenode_3_w(26);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2000w(0) <= x_prenode_3_w(27);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2008w(0) <= x_prenode_3_w(28);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2016w(0) <= x_prenode_3_w(29);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1800w(0) <= x_prenode_3_w(2);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2024w(0) <= x_prenode_3_w(30);
	wire_ccc_cordic_m_w_x_prenode_3_w_range2032w(0) <= x_prenode_3_w(31);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1808w(0) <= x_prenode_3_w(3);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1816w(0) <= x_prenode_3_w(4);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1824w(0) <= x_prenode_3_w(5);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1832w(0) <= x_prenode_3_w(6);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1840w(0) <= x_prenode_3_w(7);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1848w(0) <= x_prenode_3_w(8);
	wire_ccc_cordic_m_w_x_prenode_3_w_range1856w(0) <= x_prenode_3_w(9);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2573w(0) <= x_prenode_4_w(0);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2655w(0) <= x_prenode_4_w(10);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2663w(0) <= x_prenode_4_w(11);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2671w(0) <= x_prenode_4_w(12);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2679w(0) <= x_prenode_4_w(13);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2687w(0) <= x_prenode_4_w(14);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2695w(0) <= x_prenode_4_w(15);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2703w(0) <= x_prenode_4_w(16);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2711w(0) <= x_prenode_4_w(17);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2719w(0) <= x_prenode_4_w(18);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2727w(0) <= x_prenode_4_w(19);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2583w(0) <= x_prenode_4_w(1);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2735w(0) <= x_prenode_4_w(20);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2743w(0) <= x_prenode_4_w(21);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2751w(0) <= x_prenode_4_w(22);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2759w(0) <= x_prenode_4_w(23);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2767w(0) <= x_prenode_4_w(24);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2775w(0) <= x_prenode_4_w(25);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2783w(0) <= x_prenode_4_w(26);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2791w(0) <= x_prenode_4_w(27);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2799w(0) <= x_prenode_4_w(28);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2807w(0) <= x_prenode_4_w(29);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2591w(0) <= x_prenode_4_w(2);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2815w(0) <= x_prenode_4_w(30);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2823w(0) <= x_prenode_4_w(31);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2599w(0) <= x_prenode_4_w(3);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2607w(0) <= x_prenode_4_w(4);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2615w(0) <= x_prenode_4_w(5);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2623w(0) <= x_prenode_4_w(6);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2631w(0) <= x_prenode_4_w(7);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2639w(0) <= x_prenode_4_w(8);
	wire_ccc_cordic_m_w_x_prenode_4_w_range2647w(0) <= x_prenode_4_w(9);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3359w(0) <= x_prenode_5_w(0);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3441w(0) <= x_prenode_5_w(10);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3449w(0) <= x_prenode_5_w(11);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3457w(0) <= x_prenode_5_w(12);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3465w(0) <= x_prenode_5_w(13);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3473w(0) <= x_prenode_5_w(14);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3481w(0) <= x_prenode_5_w(15);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3489w(0) <= x_prenode_5_w(16);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3497w(0) <= x_prenode_5_w(17);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3505w(0) <= x_prenode_5_w(18);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3513w(0) <= x_prenode_5_w(19);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3369w(0) <= x_prenode_5_w(1);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3521w(0) <= x_prenode_5_w(20);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3529w(0) <= x_prenode_5_w(21);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3537w(0) <= x_prenode_5_w(22);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3545w(0) <= x_prenode_5_w(23);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3553w(0) <= x_prenode_5_w(24);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3561w(0) <= x_prenode_5_w(25);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3569w(0) <= x_prenode_5_w(26);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3577w(0) <= x_prenode_5_w(27);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3585w(0) <= x_prenode_5_w(28);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3593w(0) <= x_prenode_5_w(29);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3377w(0) <= x_prenode_5_w(2);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3601w(0) <= x_prenode_5_w(30);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3609w(0) <= x_prenode_5_w(31);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3385w(0) <= x_prenode_5_w(3);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3393w(0) <= x_prenode_5_w(4);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3401w(0) <= x_prenode_5_w(5);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3409w(0) <= x_prenode_5_w(6);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3417w(0) <= x_prenode_5_w(7);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3425w(0) <= x_prenode_5_w(8);
	wire_ccc_cordic_m_w_x_prenode_5_w_range3433w(0) <= x_prenode_5_w(9);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4140w(0) <= x_prenode_6_w(0);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4222w(0) <= x_prenode_6_w(10);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4230w(0) <= x_prenode_6_w(11);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4238w(0) <= x_prenode_6_w(12);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4246w(0) <= x_prenode_6_w(13);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4254w(0) <= x_prenode_6_w(14);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4262w(0) <= x_prenode_6_w(15);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4270w(0) <= x_prenode_6_w(16);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4278w(0) <= x_prenode_6_w(17);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4286w(0) <= x_prenode_6_w(18);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4294w(0) <= x_prenode_6_w(19);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4150w(0) <= x_prenode_6_w(1);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4302w(0) <= x_prenode_6_w(20);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4310w(0) <= x_prenode_6_w(21);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4318w(0) <= x_prenode_6_w(22);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4326w(0) <= x_prenode_6_w(23);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4334w(0) <= x_prenode_6_w(24);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4342w(0) <= x_prenode_6_w(25);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4350w(0) <= x_prenode_6_w(26);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4358w(0) <= x_prenode_6_w(27);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4366w(0) <= x_prenode_6_w(28);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4374w(0) <= x_prenode_6_w(29);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4158w(0) <= x_prenode_6_w(2);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4382w(0) <= x_prenode_6_w(30);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4390w(0) <= x_prenode_6_w(31);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4166w(0) <= x_prenode_6_w(3);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4174w(0) <= x_prenode_6_w(4);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4182w(0) <= x_prenode_6_w(5);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4190w(0) <= x_prenode_6_w(6);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4198w(0) <= x_prenode_6_w(7);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4206w(0) <= x_prenode_6_w(8);
	wire_ccc_cordic_m_w_x_prenode_6_w_range4214w(0) <= x_prenode_6_w(9);
	wire_ccc_cordic_m_w_x_prenode_7_w_range4916w(0) <= x_prenode_7_w(0);
	wire_ccc_cordic_m_w_x_prenode_7_w_range4998w(0) <= x_prenode_7_w(10);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5006w(0) <= x_prenode_7_w(11);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5014w(0) <= x_prenode_7_w(12);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5022w(0) <= x_prenode_7_w(13);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5030w(0) <= x_prenode_7_w(14);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5038w(0) <= x_prenode_7_w(15);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5046w(0) <= x_prenode_7_w(16);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5054w(0) <= x_prenode_7_w(17);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5062w(0) <= x_prenode_7_w(18);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5070w(0) <= x_prenode_7_w(19);
	wire_ccc_cordic_m_w_x_prenode_7_w_range4926w(0) <= x_prenode_7_w(1);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5078w(0) <= x_prenode_7_w(20);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5086w(0) <= x_prenode_7_w(21);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5094w(0) <= x_prenode_7_w(22);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5102w(0) <= x_prenode_7_w(23);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5110w(0) <= x_prenode_7_w(24);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5118w(0) <= x_prenode_7_w(25);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5126w(0) <= x_prenode_7_w(26);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5134w(0) <= x_prenode_7_w(27);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5142w(0) <= x_prenode_7_w(28);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5150w(0) <= x_prenode_7_w(29);
	wire_ccc_cordic_m_w_x_prenode_7_w_range4934w(0) <= x_prenode_7_w(2);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5158w(0) <= x_prenode_7_w(30);
	wire_ccc_cordic_m_w_x_prenode_7_w_range5166w(0) <= x_prenode_7_w(31);
	wire_ccc_cordic_m_w_x_prenode_7_w_range4942w(0) <= x_prenode_7_w(3);
	wire_ccc_cordic_m_w_x_prenode_7_w_range4950w(0) <= x_prenode_7_w(4);
	wire_ccc_cordic_m_w_x_prenode_7_w_range4958w(0) <= x_prenode_7_w(5);
	wire_ccc_cordic_m_w_x_prenode_7_w_range4966w(0) <= x_prenode_7_w(6);
	wire_ccc_cordic_m_w_x_prenode_7_w_range4974w(0) <= x_prenode_7_w(7);
	wire_ccc_cordic_m_w_x_prenode_7_w_range4982w(0) <= x_prenode_7_w(8);
	wire_ccc_cordic_m_w_x_prenode_7_w_range4990w(0) <= x_prenode_7_w(9);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5687w(0) <= x_prenode_8_w(0);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5769w(0) <= x_prenode_8_w(10);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5777w(0) <= x_prenode_8_w(11);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5785w(0) <= x_prenode_8_w(12);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5793w(0) <= x_prenode_8_w(13);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5801w(0) <= x_prenode_8_w(14);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5809w(0) <= x_prenode_8_w(15);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5817w(0) <= x_prenode_8_w(16);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5825w(0) <= x_prenode_8_w(17);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5833w(0) <= x_prenode_8_w(18);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5841w(0) <= x_prenode_8_w(19);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5697w(0) <= x_prenode_8_w(1);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5849w(0) <= x_prenode_8_w(20);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5857w(0) <= x_prenode_8_w(21);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5865w(0) <= x_prenode_8_w(22);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5873w(0) <= x_prenode_8_w(23);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5881w(0) <= x_prenode_8_w(24);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5889w(0) <= x_prenode_8_w(25);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5897w(0) <= x_prenode_8_w(26);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5905w(0) <= x_prenode_8_w(27);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5913w(0) <= x_prenode_8_w(28);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5921w(0) <= x_prenode_8_w(29);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5705w(0) <= x_prenode_8_w(2);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5929w(0) <= x_prenode_8_w(30);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5937w(0) <= x_prenode_8_w(31);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5713w(0) <= x_prenode_8_w(3);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5721w(0) <= x_prenode_8_w(4);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5729w(0) <= x_prenode_8_w(5);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5737w(0) <= x_prenode_8_w(6);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5745w(0) <= x_prenode_8_w(7);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5753w(0) <= x_prenode_8_w(8);
	wire_ccc_cordic_m_w_x_prenode_8_w_range5761w(0) <= x_prenode_8_w(9);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6453w(0) <= x_prenode_9_w(0);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6535w(0) <= x_prenode_9_w(10);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6543w(0) <= x_prenode_9_w(11);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6551w(0) <= x_prenode_9_w(12);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6559w(0) <= x_prenode_9_w(13);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6567w(0) <= x_prenode_9_w(14);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6575w(0) <= x_prenode_9_w(15);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6583w(0) <= x_prenode_9_w(16);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6591w(0) <= x_prenode_9_w(17);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6599w(0) <= x_prenode_9_w(18);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6607w(0) <= x_prenode_9_w(19);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6463w(0) <= x_prenode_9_w(1);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6615w(0) <= x_prenode_9_w(20);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6623w(0) <= x_prenode_9_w(21);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6631w(0) <= x_prenode_9_w(22);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6639w(0) <= x_prenode_9_w(23);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6647w(0) <= x_prenode_9_w(24);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6655w(0) <= x_prenode_9_w(25);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6663w(0) <= x_prenode_9_w(26);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6671w(0) <= x_prenode_9_w(27);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6679w(0) <= x_prenode_9_w(28);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6687w(0) <= x_prenode_9_w(29);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6471w(0) <= x_prenode_9_w(2);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6695w(0) <= x_prenode_9_w(30);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6703w(0) <= x_prenode_9_w(31);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6479w(0) <= x_prenode_9_w(3);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6487w(0) <= x_prenode_9_w(4);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6495w(0) <= x_prenode_9_w(5);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6503w(0) <= x_prenode_9_w(6);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6511w(0) <= x_prenode_9_w(7);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6519w(0) <= x_prenode_9_w(8);
	wire_ccc_cordic_m_w_x_prenode_9_w_range6527w(0) <= x_prenode_9_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7019w(0) <= x_prenodeone_10_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7078w(0) <= x_prenodeone_10_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7084w(0) <= x_prenodeone_10_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7090w(0) <= x_prenodeone_10_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7096w(0) <= x_prenodeone_10_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7102w(0) <= x_prenodeone_10_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7108w(0) <= x_prenodeone_10_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7114w(0) <= x_prenodeone_10_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7120w(0) <= x_prenodeone_10_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7126w(0) <= x_prenodeone_10_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7132w(0) <= x_prenodeone_10_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7024w(0) <= x_prenodeone_10_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7138w(0) <= x_prenodeone_10_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7144w(0) <= x_prenodeone_10_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7148w(0) <= x_prenodeone_10_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range6970w(0) <= x_prenodeone_10_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range6975w(0) <= x_prenodeone_10_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range6977w(0) <= x_prenodeone_10_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range6979w(0) <= x_prenodeone_10_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range6981w(0) <= x_prenodeone_10_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range6983w(0) <= x_prenodeone_10_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range6985w(0) <= x_prenodeone_10_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7030w(0) <= x_prenodeone_10_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range6987w(0) <= x_prenodeone_10_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range6989w(0) <= x_prenodeone_10_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7036w(0) <= x_prenodeone_10_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7042w(0) <= x_prenodeone_10_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7048w(0) <= x_prenodeone_10_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7054w(0) <= x_prenodeone_10_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7060w(0) <= x_prenodeone_10_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7066w(0) <= x_prenodeone_10_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_10_w_range7072w(0) <= x_prenodeone_10_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7784w(0) <= x_prenodeone_11_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7843w(0) <= x_prenodeone_11_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7849w(0) <= x_prenodeone_11_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7855w(0) <= x_prenodeone_11_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7861w(0) <= x_prenodeone_11_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7867w(0) <= x_prenodeone_11_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7873w(0) <= x_prenodeone_11_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7879w(0) <= x_prenodeone_11_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7885w(0) <= x_prenodeone_11_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7891w(0) <= x_prenodeone_11_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7897w(0) <= x_prenodeone_11_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7789w(0) <= x_prenodeone_11_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7903w(0) <= x_prenodeone_11_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7907w(0) <= x_prenodeone_11_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7731w(0) <= x_prenodeone_11_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7736w(0) <= x_prenodeone_11_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7738w(0) <= x_prenodeone_11_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7740w(0) <= x_prenodeone_11_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7742w(0) <= x_prenodeone_11_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7744w(0) <= x_prenodeone_11_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7746w(0) <= x_prenodeone_11_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7748w(0) <= x_prenodeone_11_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7795w(0) <= x_prenodeone_11_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7750w(0) <= x_prenodeone_11_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7752w(0) <= x_prenodeone_11_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7801w(0) <= x_prenodeone_11_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7807w(0) <= x_prenodeone_11_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7813w(0) <= x_prenodeone_11_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7819w(0) <= x_prenodeone_11_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7825w(0) <= x_prenodeone_11_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7831w(0) <= x_prenodeone_11_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_11_w_range7837w(0) <= x_prenodeone_11_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8544w(0) <= x_prenodeone_12_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8603w(0) <= x_prenodeone_12_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8609w(0) <= x_prenodeone_12_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8615w(0) <= x_prenodeone_12_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8621w(0) <= x_prenodeone_12_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8627w(0) <= x_prenodeone_12_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8633w(0) <= x_prenodeone_12_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8639w(0) <= x_prenodeone_12_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8645w(0) <= x_prenodeone_12_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8651w(0) <= x_prenodeone_12_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8657w(0) <= x_prenodeone_12_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8549w(0) <= x_prenodeone_12_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8661w(0) <= x_prenodeone_12_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8487w(0) <= x_prenodeone_12_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8492w(0) <= x_prenodeone_12_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8494w(0) <= x_prenodeone_12_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8496w(0) <= x_prenodeone_12_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8498w(0) <= x_prenodeone_12_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8500w(0) <= x_prenodeone_12_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8502w(0) <= x_prenodeone_12_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8504w(0) <= x_prenodeone_12_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8506w(0) <= x_prenodeone_12_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8555w(0) <= x_prenodeone_12_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8508w(0) <= x_prenodeone_12_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8510w(0) <= x_prenodeone_12_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8561w(0) <= x_prenodeone_12_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8567w(0) <= x_prenodeone_12_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8573w(0) <= x_prenodeone_12_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8579w(0) <= x_prenodeone_12_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8585w(0) <= x_prenodeone_12_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8591w(0) <= x_prenodeone_12_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_12_w_range8597w(0) <= x_prenodeone_12_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9299w(0) <= x_prenodeone_13_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9358w(0) <= x_prenodeone_13_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9364w(0) <= x_prenodeone_13_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9370w(0) <= x_prenodeone_13_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9376w(0) <= x_prenodeone_13_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9382w(0) <= x_prenodeone_13_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9388w(0) <= x_prenodeone_13_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9394w(0) <= x_prenodeone_13_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9400w(0) <= x_prenodeone_13_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9406w(0) <= x_prenodeone_13_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9410w(0) <= x_prenodeone_13_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9304w(0) <= x_prenodeone_13_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9238w(0) <= x_prenodeone_13_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9243w(0) <= x_prenodeone_13_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9245w(0) <= x_prenodeone_13_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9247w(0) <= x_prenodeone_13_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9249w(0) <= x_prenodeone_13_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9251w(0) <= x_prenodeone_13_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9253w(0) <= x_prenodeone_13_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9255w(0) <= x_prenodeone_13_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9257w(0) <= x_prenodeone_13_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9259w(0) <= x_prenodeone_13_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9310w(0) <= x_prenodeone_13_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9261w(0) <= x_prenodeone_13_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9263w(0) <= x_prenodeone_13_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9316w(0) <= x_prenodeone_13_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9322w(0) <= x_prenodeone_13_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9328w(0) <= x_prenodeone_13_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9334w(0) <= x_prenodeone_13_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9340w(0) <= x_prenodeone_13_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9346w(0) <= x_prenodeone_13_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_13_w_range9352w(0) <= x_prenodeone_13_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range719w(0) <= x_prenodeone_2_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range778w(0) <= x_prenodeone_2_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range784w(0) <= x_prenodeone_2_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range790w(0) <= x_prenodeone_2_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range796w(0) <= x_prenodeone_2_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range802w(0) <= x_prenodeone_2_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range808w(0) <= x_prenodeone_2_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range814w(0) <= x_prenodeone_2_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range820w(0) <= x_prenodeone_2_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range826w(0) <= x_prenodeone_2_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range832w(0) <= x_prenodeone_2_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range724w(0) <= x_prenodeone_2_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range838w(0) <= x_prenodeone_2_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range844w(0) <= x_prenodeone_2_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range850w(0) <= x_prenodeone_2_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range856w(0) <= x_prenodeone_2_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range862w(0) <= x_prenodeone_2_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range868w(0) <= x_prenodeone_2_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range874w(0) <= x_prenodeone_2_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range880w(0) <= x_prenodeone_2_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range886w(0) <= x_prenodeone_2_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range892w(0) <= x_prenodeone_2_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range730w(0) <= x_prenodeone_2_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range896w(0) <= x_prenodeone_2_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range702w(0) <= x_prenodeone_2_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range736w(0) <= x_prenodeone_2_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range742w(0) <= x_prenodeone_2_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range748w(0) <= x_prenodeone_2_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range754w(0) <= x_prenodeone_2_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range760w(0) <= x_prenodeone_2_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range766w(0) <= x_prenodeone_2_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_2_w_range772w(0) <= x_prenodeone_2_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1524w(0) <= x_prenodeone_3_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1583w(0) <= x_prenodeone_3_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1589w(0) <= x_prenodeone_3_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1595w(0) <= x_prenodeone_3_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1601w(0) <= x_prenodeone_3_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1607w(0) <= x_prenodeone_3_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1613w(0) <= x_prenodeone_3_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1619w(0) <= x_prenodeone_3_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1625w(0) <= x_prenodeone_3_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1631w(0) <= x_prenodeone_3_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1637w(0) <= x_prenodeone_3_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1529w(0) <= x_prenodeone_3_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1643w(0) <= x_prenodeone_3_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1649w(0) <= x_prenodeone_3_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1655w(0) <= x_prenodeone_3_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1661w(0) <= x_prenodeone_3_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1667w(0) <= x_prenodeone_3_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1673w(0) <= x_prenodeone_3_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1679w(0) <= x_prenodeone_3_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1685w(0) <= x_prenodeone_3_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1691w(0) <= x_prenodeone_3_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1695w(0) <= x_prenodeone_3_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1535w(0) <= x_prenodeone_3_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1503w(0) <= x_prenodeone_3_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1508w(0) <= x_prenodeone_3_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1541w(0) <= x_prenodeone_3_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1547w(0) <= x_prenodeone_3_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1553w(0) <= x_prenodeone_3_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1559w(0) <= x_prenodeone_3_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1565w(0) <= x_prenodeone_3_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1571w(0) <= x_prenodeone_3_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_3_w_range1577w(0) <= x_prenodeone_3_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2324w(0) <= x_prenodeone_4_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2383w(0) <= x_prenodeone_4_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2389w(0) <= x_prenodeone_4_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2395w(0) <= x_prenodeone_4_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2401w(0) <= x_prenodeone_4_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2407w(0) <= x_prenodeone_4_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2413w(0) <= x_prenodeone_4_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2419w(0) <= x_prenodeone_4_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2425w(0) <= x_prenodeone_4_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2431w(0) <= x_prenodeone_4_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2437w(0) <= x_prenodeone_4_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2329w(0) <= x_prenodeone_4_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2443w(0) <= x_prenodeone_4_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2449w(0) <= x_prenodeone_4_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2455w(0) <= x_prenodeone_4_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2461w(0) <= x_prenodeone_4_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2467w(0) <= x_prenodeone_4_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2473w(0) <= x_prenodeone_4_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2479w(0) <= x_prenodeone_4_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2485w(0) <= x_prenodeone_4_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2489w(0) <= x_prenodeone_4_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2299w(0) <= x_prenodeone_4_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2335w(0) <= x_prenodeone_4_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2304w(0) <= x_prenodeone_4_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2306w(0) <= x_prenodeone_4_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2341w(0) <= x_prenodeone_4_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2347w(0) <= x_prenodeone_4_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2353w(0) <= x_prenodeone_4_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2359w(0) <= x_prenodeone_4_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2365w(0) <= x_prenodeone_4_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2371w(0) <= x_prenodeone_4_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_4_w_range2377w(0) <= x_prenodeone_4_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3119w(0) <= x_prenodeone_5_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3178w(0) <= x_prenodeone_5_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3184w(0) <= x_prenodeone_5_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3190w(0) <= x_prenodeone_5_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3196w(0) <= x_prenodeone_5_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3202w(0) <= x_prenodeone_5_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3208w(0) <= x_prenodeone_5_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3214w(0) <= x_prenodeone_5_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3220w(0) <= x_prenodeone_5_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3226w(0) <= x_prenodeone_5_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3232w(0) <= x_prenodeone_5_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3124w(0) <= x_prenodeone_5_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3238w(0) <= x_prenodeone_5_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3244w(0) <= x_prenodeone_5_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3250w(0) <= x_prenodeone_5_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3256w(0) <= x_prenodeone_5_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3262w(0) <= x_prenodeone_5_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3268w(0) <= x_prenodeone_5_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3274w(0) <= x_prenodeone_5_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3278w(0) <= x_prenodeone_5_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3090w(0) <= x_prenodeone_5_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3095w(0) <= x_prenodeone_5_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3130w(0) <= x_prenodeone_5_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3097w(0) <= x_prenodeone_5_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3099w(0) <= x_prenodeone_5_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3136w(0) <= x_prenodeone_5_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3142w(0) <= x_prenodeone_5_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3148w(0) <= x_prenodeone_5_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3154w(0) <= x_prenodeone_5_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3160w(0) <= x_prenodeone_5_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3166w(0) <= x_prenodeone_5_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_5_w_range3172w(0) <= x_prenodeone_5_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3909w(0) <= x_prenodeone_6_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3968w(0) <= x_prenodeone_6_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3974w(0) <= x_prenodeone_6_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3980w(0) <= x_prenodeone_6_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3986w(0) <= x_prenodeone_6_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3992w(0) <= x_prenodeone_6_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3998w(0) <= x_prenodeone_6_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4004w(0) <= x_prenodeone_6_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4010w(0) <= x_prenodeone_6_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4016w(0) <= x_prenodeone_6_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4022w(0) <= x_prenodeone_6_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3914w(0) <= x_prenodeone_6_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4028w(0) <= x_prenodeone_6_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4034w(0) <= x_prenodeone_6_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4040w(0) <= x_prenodeone_6_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4046w(0) <= x_prenodeone_6_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4052w(0) <= x_prenodeone_6_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4058w(0) <= x_prenodeone_6_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range4062w(0) <= x_prenodeone_6_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3876w(0) <= x_prenodeone_6_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3881w(0) <= x_prenodeone_6_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3883w(0) <= x_prenodeone_6_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3920w(0) <= x_prenodeone_6_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3885w(0) <= x_prenodeone_6_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3887w(0) <= x_prenodeone_6_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3926w(0) <= x_prenodeone_6_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3932w(0) <= x_prenodeone_6_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3938w(0) <= x_prenodeone_6_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3944w(0) <= x_prenodeone_6_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3950w(0) <= x_prenodeone_6_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3956w(0) <= x_prenodeone_6_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_6_w_range3962w(0) <= x_prenodeone_6_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4694w(0) <= x_prenodeone_7_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4753w(0) <= x_prenodeone_7_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4759w(0) <= x_prenodeone_7_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4765w(0) <= x_prenodeone_7_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4771w(0) <= x_prenodeone_7_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4777w(0) <= x_prenodeone_7_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4783w(0) <= x_prenodeone_7_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4789w(0) <= x_prenodeone_7_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4795w(0) <= x_prenodeone_7_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4801w(0) <= x_prenodeone_7_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4807w(0) <= x_prenodeone_7_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4699w(0) <= x_prenodeone_7_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4813w(0) <= x_prenodeone_7_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4819w(0) <= x_prenodeone_7_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4825w(0) <= x_prenodeone_7_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4831w(0) <= x_prenodeone_7_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4837w(0) <= x_prenodeone_7_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4841w(0) <= x_prenodeone_7_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4657w(0) <= x_prenodeone_7_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4662w(0) <= x_prenodeone_7_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4664w(0) <= x_prenodeone_7_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4666w(0) <= x_prenodeone_7_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4705w(0) <= x_prenodeone_7_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4668w(0) <= x_prenodeone_7_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4670w(0) <= x_prenodeone_7_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4711w(0) <= x_prenodeone_7_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4717w(0) <= x_prenodeone_7_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4723w(0) <= x_prenodeone_7_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4729w(0) <= x_prenodeone_7_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4735w(0) <= x_prenodeone_7_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4741w(0) <= x_prenodeone_7_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_7_w_range4747w(0) <= x_prenodeone_7_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5474w(0) <= x_prenodeone_8_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5533w(0) <= x_prenodeone_8_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5539w(0) <= x_prenodeone_8_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5545w(0) <= x_prenodeone_8_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5551w(0) <= x_prenodeone_8_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5557w(0) <= x_prenodeone_8_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5563w(0) <= x_prenodeone_8_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5569w(0) <= x_prenodeone_8_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5575w(0) <= x_prenodeone_8_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5581w(0) <= x_prenodeone_8_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5587w(0) <= x_prenodeone_8_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5479w(0) <= x_prenodeone_8_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5593w(0) <= x_prenodeone_8_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5599w(0) <= x_prenodeone_8_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5605w(0) <= x_prenodeone_8_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5611w(0) <= x_prenodeone_8_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5615w(0) <= x_prenodeone_8_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5433w(0) <= x_prenodeone_8_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5438w(0) <= x_prenodeone_8_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5440w(0) <= x_prenodeone_8_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5442w(0) <= x_prenodeone_8_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5444w(0) <= x_prenodeone_8_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5485w(0) <= x_prenodeone_8_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5446w(0) <= x_prenodeone_8_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5448w(0) <= x_prenodeone_8_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5491w(0) <= x_prenodeone_8_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5497w(0) <= x_prenodeone_8_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5503w(0) <= x_prenodeone_8_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5509w(0) <= x_prenodeone_8_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5515w(0) <= x_prenodeone_8_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5521w(0) <= x_prenodeone_8_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_8_w_range5527w(0) <= x_prenodeone_8_w(9);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6249w(0) <= x_prenodeone_9_w(0);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6308w(0) <= x_prenodeone_9_w(10);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6314w(0) <= x_prenodeone_9_w(11);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6320w(0) <= x_prenodeone_9_w(12);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6326w(0) <= x_prenodeone_9_w(13);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6332w(0) <= x_prenodeone_9_w(14);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6338w(0) <= x_prenodeone_9_w(15);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6344w(0) <= x_prenodeone_9_w(16);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6350w(0) <= x_prenodeone_9_w(17);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6356w(0) <= x_prenodeone_9_w(18);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6362w(0) <= x_prenodeone_9_w(19);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6254w(0) <= x_prenodeone_9_w(1);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6368w(0) <= x_prenodeone_9_w(20);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6374w(0) <= x_prenodeone_9_w(21);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6380w(0) <= x_prenodeone_9_w(22);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6384w(0) <= x_prenodeone_9_w(23);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6204w(0) <= x_prenodeone_9_w(24);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6209w(0) <= x_prenodeone_9_w(25);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6211w(0) <= x_prenodeone_9_w(26);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6213w(0) <= x_prenodeone_9_w(27);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6215w(0) <= x_prenodeone_9_w(28);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6217w(0) <= x_prenodeone_9_w(29);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6260w(0) <= x_prenodeone_9_w(2);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6219w(0) <= x_prenodeone_9_w(30);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6221w(0) <= x_prenodeone_9_w(31);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6266w(0) <= x_prenodeone_9_w(3);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6272w(0) <= x_prenodeone_9_w(4);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6278w(0) <= x_prenodeone_9_w(5);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6284w(0) <= x_prenodeone_9_w(6);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6290w(0) <= x_prenodeone_9_w(7);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6296w(0) <= x_prenodeone_9_w(8);
	wire_ccc_cordic_m_w_x_prenodeone_9_w_range6302w(0) <= x_prenodeone_9_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7151w(0) <= x_prenodetwo_10_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7180w(0) <= x_prenodetwo_10_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7183w(0) <= x_prenodetwo_10_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7186w(0) <= x_prenodetwo_10_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7189w(0) <= x_prenodetwo_10_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7192w(0) <= x_prenodetwo_10_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7195w(0) <= x_prenodetwo_10_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7198w(0) <= x_prenodetwo_10_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7201w(0) <= x_prenodetwo_10_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7204w(0) <= x_prenodetwo_10_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7207w(0) <= x_prenodetwo_10_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7153w(0) <= x_prenodetwo_10_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range6991w(0) <= x_prenodetwo_10_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range6995w(0) <= x_prenodetwo_10_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range6997w(0) <= x_prenodetwo_10_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range6999w(0) <= x_prenodetwo_10_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7001w(0) <= x_prenodetwo_10_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7003w(0) <= x_prenodetwo_10_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7005w(0) <= x_prenodetwo_10_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7007w(0) <= x_prenodetwo_10_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7009w(0) <= x_prenodetwo_10_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7011w(0) <= x_prenodetwo_10_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7156w(0) <= x_prenodetwo_10_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7013w(0) <= x_prenodetwo_10_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7015w(0) <= x_prenodetwo_10_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7159w(0) <= x_prenodetwo_10_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7162w(0) <= x_prenodetwo_10_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7165w(0) <= x_prenodetwo_10_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7168w(0) <= x_prenodetwo_10_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7171w(0) <= x_prenodetwo_10_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7174w(0) <= x_prenodetwo_10_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_10_w_range7177w(0) <= x_prenodetwo_10_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7910w(0) <= x_prenodetwo_11_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7939w(0) <= x_prenodetwo_11_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7942w(0) <= x_prenodetwo_11_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7945w(0) <= x_prenodetwo_11_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7948w(0) <= x_prenodetwo_11_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7951w(0) <= x_prenodetwo_11_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7954w(0) <= x_prenodetwo_11_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7957w(0) <= x_prenodetwo_11_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7960w(0) <= x_prenodetwo_11_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7963w(0) <= x_prenodetwo_11_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7754w(0) <= x_prenodetwo_11_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7912w(0) <= x_prenodetwo_11_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7758w(0) <= x_prenodetwo_11_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7760w(0) <= x_prenodetwo_11_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7762w(0) <= x_prenodetwo_11_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7764w(0) <= x_prenodetwo_11_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7766w(0) <= x_prenodetwo_11_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7768w(0) <= x_prenodetwo_11_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7770w(0) <= x_prenodetwo_11_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7772w(0) <= x_prenodetwo_11_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7774w(0) <= x_prenodetwo_11_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7776w(0) <= x_prenodetwo_11_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7915w(0) <= x_prenodetwo_11_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7778w(0) <= x_prenodetwo_11_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7780w(0) <= x_prenodetwo_11_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7918w(0) <= x_prenodetwo_11_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7921w(0) <= x_prenodetwo_11_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7924w(0) <= x_prenodetwo_11_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7927w(0) <= x_prenodetwo_11_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7930w(0) <= x_prenodetwo_11_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7933w(0) <= x_prenodetwo_11_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_11_w_range7936w(0) <= x_prenodetwo_11_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8664w(0) <= x_prenodetwo_12_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8693w(0) <= x_prenodetwo_12_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8696w(0) <= x_prenodetwo_12_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8699w(0) <= x_prenodetwo_12_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8702w(0) <= x_prenodetwo_12_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8705w(0) <= x_prenodetwo_12_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8708w(0) <= x_prenodetwo_12_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8711w(0) <= x_prenodetwo_12_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8714w(0) <= x_prenodetwo_12_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8512w(0) <= x_prenodetwo_12_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8516w(0) <= x_prenodetwo_12_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8666w(0) <= x_prenodetwo_12_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8518w(0) <= x_prenodetwo_12_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8520w(0) <= x_prenodetwo_12_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8522w(0) <= x_prenodetwo_12_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8524w(0) <= x_prenodetwo_12_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8526w(0) <= x_prenodetwo_12_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8528w(0) <= x_prenodetwo_12_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8530w(0) <= x_prenodetwo_12_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8532w(0) <= x_prenodetwo_12_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8534w(0) <= x_prenodetwo_12_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8536w(0) <= x_prenodetwo_12_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8669w(0) <= x_prenodetwo_12_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8538w(0) <= x_prenodetwo_12_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8540w(0) <= x_prenodetwo_12_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8672w(0) <= x_prenodetwo_12_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8675w(0) <= x_prenodetwo_12_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8678w(0) <= x_prenodetwo_12_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8681w(0) <= x_prenodetwo_12_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8684w(0) <= x_prenodetwo_12_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8687w(0) <= x_prenodetwo_12_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_12_w_range8690w(0) <= x_prenodetwo_12_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9413w(0) <= x_prenodetwo_13_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9442w(0) <= x_prenodetwo_13_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9445w(0) <= x_prenodetwo_13_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9448w(0) <= x_prenodetwo_13_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9451w(0) <= x_prenodetwo_13_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9454w(0) <= x_prenodetwo_13_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9457w(0) <= x_prenodetwo_13_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9460w(0) <= x_prenodetwo_13_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9265w(0) <= x_prenodetwo_13_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9269w(0) <= x_prenodetwo_13_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9271w(0) <= x_prenodetwo_13_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9415w(0) <= x_prenodetwo_13_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9273w(0) <= x_prenodetwo_13_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9275w(0) <= x_prenodetwo_13_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9277w(0) <= x_prenodetwo_13_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9279w(0) <= x_prenodetwo_13_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9281w(0) <= x_prenodetwo_13_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9283w(0) <= x_prenodetwo_13_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9285w(0) <= x_prenodetwo_13_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9287w(0) <= x_prenodetwo_13_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9289w(0) <= x_prenodetwo_13_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9291w(0) <= x_prenodetwo_13_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9418w(0) <= x_prenodetwo_13_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9293w(0) <= x_prenodetwo_13_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9295w(0) <= x_prenodetwo_13_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9421w(0) <= x_prenodetwo_13_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9424w(0) <= x_prenodetwo_13_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9427w(0) <= x_prenodetwo_13_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9430w(0) <= x_prenodetwo_13_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9433w(0) <= x_prenodetwo_13_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9436w(0) <= x_prenodetwo_13_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_13_w_range9439w(0) <= x_prenodetwo_13_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range899w(0) <= x_prenodetwo_2_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range928w(0) <= x_prenodetwo_2_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range931w(0) <= x_prenodetwo_2_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range934w(0) <= x_prenodetwo_2_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range937w(0) <= x_prenodetwo_2_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range940w(0) <= x_prenodetwo_2_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range943w(0) <= x_prenodetwo_2_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range946w(0) <= x_prenodetwo_2_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range949w(0) <= x_prenodetwo_2_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range952w(0) <= x_prenodetwo_2_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range955w(0) <= x_prenodetwo_2_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range901w(0) <= x_prenodetwo_2_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range958w(0) <= x_prenodetwo_2_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range961w(0) <= x_prenodetwo_2_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range964w(0) <= x_prenodetwo_2_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range967w(0) <= x_prenodetwo_2_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range970w(0) <= x_prenodetwo_2_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range973w(0) <= x_prenodetwo_2_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range976w(0) <= x_prenodetwo_2_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range979w(0) <= x_prenodetwo_2_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range707w(0) <= x_prenodetwo_2_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range711w(0) <= x_prenodetwo_2_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range904w(0) <= x_prenodetwo_2_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range713w(0) <= x_prenodetwo_2_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range715w(0) <= x_prenodetwo_2_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range907w(0) <= x_prenodetwo_2_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range910w(0) <= x_prenodetwo_2_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range913w(0) <= x_prenodetwo_2_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range916w(0) <= x_prenodetwo_2_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range919w(0) <= x_prenodetwo_2_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range922w(0) <= x_prenodetwo_2_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_2_w_range925w(0) <= x_prenodetwo_2_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1698w(0) <= x_prenodetwo_3_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1727w(0) <= x_prenodetwo_3_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1730w(0) <= x_prenodetwo_3_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1733w(0) <= x_prenodetwo_3_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1736w(0) <= x_prenodetwo_3_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1739w(0) <= x_prenodetwo_3_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1742w(0) <= x_prenodetwo_3_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1745w(0) <= x_prenodetwo_3_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1748w(0) <= x_prenodetwo_3_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1751w(0) <= x_prenodetwo_3_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1754w(0) <= x_prenodetwo_3_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1700w(0) <= x_prenodetwo_3_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1757w(0) <= x_prenodetwo_3_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1760w(0) <= x_prenodetwo_3_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1763w(0) <= x_prenodetwo_3_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1766w(0) <= x_prenodetwo_3_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1769w(0) <= x_prenodetwo_3_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1772w(0) <= x_prenodetwo_3_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1775w(0) <= x_prenodetwo_3_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1510w(0) <= x_prenodetwo_3_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1514w(0) <= x_prenodetwo_3_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1516w(0) <= x_prenodetwo_3_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1703w(0) <= x_prenodetwo_3_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1518w(0) <= x_prenodetwo_3_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1520w(0) <= x_prenodetwo_3_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1706w(0) <= x_prenodetwo_3_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1709w(0) <= x_prenodetwo_3_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1712w(0) <= x_prenodetwo_3_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1715w(0) <= x_prenodetwo_3_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1718w(0) <= x_prenodetwo_3_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1721w(0) <= x_prenodetwo_3_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_3_w_range1724w(0) <= x_prenodetwo_3_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2492w(0) <= x_prenodetwo_4_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2521w(0) <= x_prenodetwo_4_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2524w(0) <= x_prenodetwo_4_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2527w(0) <= x_prenodetwo_4_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2530w(0) <= x_prenodetwo_4_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2533w(0) <= x_prenodetwo_4_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2536w(0) <= x_prenodetwo_4_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2539w(0) <= x_prenodetwo_4_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2542w(0) <= x_prenodetwo_4_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2545w(0) <= x_prenodetwo_4_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2548w(0) <= x_prenodetwo_4_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2494w(0) <= x_prenodetwo_4_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2551w(0) <= x_prenodetwo_4_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2554w(0) <= x_prenodetwo_4_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2557w(0) <= x_prenodetwo_4_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2560w(0) <= x_prenodetwo_4_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2563w(0) <= x_prenodetwo_4_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2566w(0) <= x_prenodetwo_4_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2308w(0) <= x_prenodetwo_4_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2312w(0) <= x_prenodetwo_4_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2314w(0) <= x_prenodetwo_4_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2316w(0) <= x_prenodetwo_4_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2497w(0) <= x_prenodetwo_4_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2318w(0) <= x_prenodetwo_4_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2320w(0) <= x_prenodetwo_4_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2500w(0) <= x_prenodetwo_4_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2503w(0) <= x_prenodetwo_4_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2506w(0) <= x_prenodetwo_4_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2509w(0) <= x_prenodetwo_4_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2512w(0) <= x_prenodetwo_4_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2515w(0) <= x_prenodetwo_4_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_4_w_range2518w(0) <= x_prenodetwo_4_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3281w(0) <= x_prenodetwo_5_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3310w(0) <= x_prenodetwo_5_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3313w(0) <= x_prenodetwo_5_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3316w(0) <= x_prenodetwo_5_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3319w(0) <= x_prenodetwo_5_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3322w(0) <= x_prenodetwo_5_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3325w(0) <= x_prenodetwo_5_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3328w(0) <= x_prenodetwo_5_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3331w(0) <= x_prenodetwo_5_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3334w(0) <= x_prenodetwo_5_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3337w(0) <= x_prenodetwo_5_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3283w(0) <= x_prenodetwo_5_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3340w(0) <= x_prenodetwo_5_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3343w(0) <= x_prenodetwo_5_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3346w(0) <= x_prenodetwo_5_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3349w(0) <= x_prenodetwo_5_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3352w(0) <= x_prenodetwo_5_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3101w(0) <= x_prenodetwo_5_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3105w(0) <= x_prenodetwo_5_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3107w(0) <= x_prenodetwo_5_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3109w(0) <= x_prenodetwo_5_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3111w(0) <= x_prenodetwo_5_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3286w(0) <= x_prenodetwo_5_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3113w(0) <= x_prenodetwo_5_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3115w(0) <= x_prenodetwo_5_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3289w(0) <= x_prenodetwo_5_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3292w(0) <= x_prenodetwo_5_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3295w(0) <= x_prenodetwo_5_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3298w(0) <= x_prenodetwo_5_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3301w(0) <= x_prenodetwo_5_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3304w(0) <= x_prenodetwo_5_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_5_w_range3307w(0) <= x_prenodetwo_5_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4065w(0) <= x_prenodetwo_6_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4094w(0) <= x_prenodetwo_6_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4097w(0) <= x_prenodetwo_6_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4100w(0) <= x_prenodetwo_6_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4103w(0) <= x_prenodetwo_6_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4106w(0) <= x_prenodetwo_6_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4109w(0) <= x_prenodetwo_6_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4112w(0) <= x_prenodetwo_6_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4115w(0) <= x_prenodetwo_6_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4118w(0) <= x_prenodetwo_6_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4121w(0) <= x_prenodetwo_6_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4067w(0) <= x_prenodetwo_6_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4124w(0) <= x_prenodetwo_6_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4127w(0) <= x_prenodetwo_6_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4130w(0) <= x_prenodetwo_6_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4133w(0) <= x_prenodetwo_6_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3889w(0) <= x_prenodetwo_6_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3893w(0) <= x_prenodetwo_6_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3895w(0) <= x_prenodetwo_6_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3897w(0) <= x_prenodetwo_6_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3899w(0) <= x_prenodetwo_6_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3901w(0) <= x_prenodetwo_6_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4070w(0) <= x_prenodetwo_6_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3903w(0) <= x_prenodetwo_6_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range3905w(0) <= x_prenodetwo_6_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4073w(0) <= x_prenodetwo_6_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4076w(0) <= x_prenodetwo_6_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4079w(0) <= x_prenodetwo_6_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4082w(0) <= x_prenodetwo_6_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4085w(0) <= x_prenodetwo_6_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4088w(0) <= x_prenodetwo_6_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_6_w_range4091w(0) <= x_prenodetwo_6_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4844w(0) <= x_prenodetwo_7_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4873w(0) <= x_prenodetwo_7_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4876w(0) <= x_prenodetwo_7_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4879w(0) <= x_prenodetwo_7_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4882w(0) <= x_prenodetwo_7_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4885w(0) <= x_prenodetwo_7_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4888w(0) <= x_prenodetwo_7_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4891w(0) <= x_prenodetwo_7_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4894w(0) <= x_prenodetwo_7_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4897w(0) <= x_prenodetwo_7_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4900w(0) <= x_prenodetwo_7_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4846w(0) <= x_prenodetwo_7_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4903w(0) <= x_prenodetwo_7_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4906w(0) <= x_prenodetwo_7_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4909w(0) <= x_prenodetwo_7_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4672w(0) <= x_prenodetwo_7_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4676w(0) <= x_prenodetwo_7_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4678w(0) <= x_prenodetwo_7_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4680w(0) <= x_prenodetwo_7_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4682w(0) <= x_prenodetwo_7_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4684w(0) <= x_prenodetwo_7_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4686w(0) <= x_prenodetwo_7_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4849w(0) <= x_prenodetwo_7_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4688w(0) <= x_prenodetwo_7_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4690w(0) <= x_prenodetwo_7_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4852w(0) <= x_prenodetwo_7_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4855w(0) <= x_prenodetwo_7_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4858w(0) <= x_prenodetwo_7_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4861w(0) <= x_prenodetwo_7_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4864w(0) <= x_prenodetwo_7_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4867w(0) <= x_prenodetwo_7_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_7_w_range4870w(0) <= x_prenodetwo_7_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5618w(0) <= x_prenodetwo_8_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5647w(0) <= x_prenodetwo_8_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5650w(0) <= x_prenodetwo_8_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5653w(0) <= x_prenodetwo_8_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5656w(0) <= x_prenodetwo_8_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5659w(0) <= x_prenodetwo_8_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5662w(0) <= x_prenodetwo_8_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5665w(0) <= x_prenodetwo_8_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5668w(0) <= x_prenodetwo_8_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5671w(0) <= x_prenodetwo_8_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5674w(0) <= x_prenodetwo_8_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5620w(0) <= x_prenodetwo_8_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5677w(0) <= x_prenodetwo_8_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5680w(0) <= x_prenodetwo_8_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5450w(0) <= x_prenodetwo_8_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5454w(0) <= x_prenodetwo_8_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5456w(0) <= x_prenodetwo_8_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5458w(0) <= x_prenodetwo_8_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5460w(0) <= x_prenodetwo_8_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5462w(0) <= x_prenodetwo_8_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5464w(0) <= x_prenodetwo_8_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5466w(0) <= x_prenodetwo_8_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5623w(0) <= x_prenodetwo_8_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5468w(0) <= x_prenodetwo_8_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5470w(0) <= x_prenodetwo_8_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5626w(0) <= x_prenodetwo_8_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5629w(0) <= x_prenodetwo_8_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5632w(0) <= x_prenodetwo_8_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5635w(0) <= x_prenodetwo_8_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5638w(0) <= x_prenodetwo_8_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5641w(0) <= x_prenodetwo_8_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_8_w_range5644w(0) <= x_prenodetwo_8_w(9);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6387w(0) <= x_prenodetwo_9_w(0);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6416w(0) <= x_prenodetwo_9_w(10);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6419w(0) <= x_prenodetwo_9_w(11);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6422w(0) <= x_prenodetwo_9_w(12);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6425w(0) <= x_prenodetwo_9_w(13);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6428w(0) <= x_prenodetwo_9_w(14);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6431w(0) <= x_prenodetwo_9_w(15);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6434w(0) <= x_prenodetwo_9_w(16);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6437w(0) <= x_prenodetwo_9_w(17);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6440w(0) <= x_prenodetwo_9_w(18);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6443w(0) <= x_prenodetwo_9_w(19);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6389w(0) <= x_prenodetwo_9_w(1);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6446w(0) <= x_prenodetwo_9_w(20);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6223w(0) <= x_prenodetwo_9_w(21);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6227w(0) <= x_prenodetwo_9_w(22);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6229w(0) <= x_prenodetwo_9_w(23);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6231w(0) <= x_prenodetwo_9_w(24);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6233w(0) <= x_prenodetwo_9_w(25);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6235w(0) <= x_prenodetwo_9_w(26);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6237w(0) <= x_prenodetwo_9_w(27);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6239w(0) <= x_prenodetwo_9_w(28);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6241w(0) <= x_prenodetwo_9_w(29);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6392w(0) <= x_prenodetwo_9_w(2);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6243w(0) <= x_prenodetwo_9_w(30);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6245w(0) <= x_prenodetwo_9_w(31);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6395w(0) <= x_prenodetwo_9_w(3);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6398w(0) <= x_prenodetwo_9_w(4);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6401w(0) <= x_prenodetwo_9_w(5);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6404w(0) <= x_prenodetwo_9_w(6);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6407w(0) <= x_prenodetwo_9_w(7);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6410w(0) <= x_prenodetwo_9_w(8);
	wire_ccc_cordic_m_w_x_prenodetwo_9_w_range6413w(0) <= x_prenodetwo_9_w(9);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7219w(0) <= y_prenode_10_w(0);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7300w(0) <= y_prenode_10_w(10);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7308w(0) <= y_prenode_10_w(11);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7316w(0) <= y_prenode_10_w(12);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7324w(0) <= y_prenode_10_w(13);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7332w(0) <= y_prenode_10_w(14);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7340w(0) <= y_prenode_10_w(15);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7348w(0) <= y_prenode_10_w(16);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7356w(0) <= y_prenode_10_w(17);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7364w(0) <= y_prenode_10_w(18);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7372w(0) <= y_prenode_10_w(19);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7228w(0) <= y_prenode_10_w(1);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7380w(0) <= y_prenode_10_w(20);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7388w(0) <= y_prenode_10_w(21);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7396w(0) <= y_prenode_10_w(22);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7404w(0) <= y_prenode_10_w(23);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7412w(0) <= y_prenode_10_w(24);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7420w(0) <= y_prenode_10_w(25);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7428w(0) <= y_prenode_10_w(26);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7436w(0) <= y_prenode_10_w(27);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7444w(0) <= y_prenode_10_w(28);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7452w(0) <= y_prenode_10_w(29);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7236w(0) <= y_prenode_10_w(2);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7460w(0) <= y_prenode_10_w(30);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7468w(0) <= y_prenode_10_w(31);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7244w(0) <= y_prenode_10_w(3);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7252w(0) <= y_prenode_10_w(4);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7260w(0) <= y_prenode_10_w(5);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7268w(0) <= y_prenode_10_w(6);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7276w(0) <= y_prenode_10_w(7);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7284w(0) <= y_prenode_10_w(8);
	wire_ccc_cordic_m_w_y_prenode_10_w_range7292w(0) <= y_prenode_10_w(9);
	wire_ccc_cordic_m_w_y_prenode_11_w_range7975w(0) <= y_prenode_11_w(0);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8056w(0) <= y_prenode_11_w(10);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8064w(0) <= y_prenode_11_w(11);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8072w(0) <= y_prenode_11_w(12);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8080w(0) <= y_prenode_11_w(13);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8088w(0) <= y_prenode_11_w(14);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8096w(0) <= y_prenode_11_w(15);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8104w(0) <= y_prenode_11_w(16);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8112w(0) <= y_prenode_11_w(17);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8120w(0) <= y_prenode_11_w(18);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8128w(0) <= y_prenode_11_w(19);
	wire_ccc_cordic_m_w_y_prenode_11_w_range7984w(0) <= y_prenode_11_w(1);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8136w(0) <= y_prenode_11_w(20);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8144w(0) <= y_prenode_11_w(21);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8152w(0) <= y_prenode_11_w(22);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8160w(0) <= y_prenode_11_w(23);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8168w(0) <= y_prenode_11_w(24);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8176w(0) <= y_prenode_11_w(25);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8184w(0) <= y_prenode_11_w(26);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8192w(0) <= y_prenode_11_w(27);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8200w(0) <= y_prenode_11_w(28);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8208w(0) <= y_prenode_11_w(29);
	wire_ccc_cordic_m_w_y_prenode_11_w_range7992w(0) <= y_prenode_11_w(2);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8216w(0) <= y_prenode_11_w(30);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8224w(0) <= y_prenode_11_w(31);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8000w(0) <= y_prenode_11_w(3);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8008w(0) <= y_prenode_11_w(4);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8016w(0) <= y_prenode_11_w(5);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8024w(0) <= y_prenode_11_w(6);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8032w(0) <= y_prenode_11_w(7);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8040w(0) <= y_prenode_11_w(8);
	wire_ccc_cordic_m_w_y_prenode_11_w_range8048w(0) <= y_prenode_11_w(9);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8726w(0) <= y_prenode_12_w(0);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8807w(0) <= y_prenode_12_w(10);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8815w(0) <= y_prenode_12_w(11);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8823w(0) <= y_prenode_12_w(12);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8831w(0) <= y_prenode_12_w(13);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8839w(0) <= y_prenode_12_w(14);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8847w(0) <= y_prenode_12_w(15);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8855w(0) <= y_prenode_12_w(16);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8863w(0) <= y_prenode_12_w(17);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8871w(0) <= y_prenode_12_w(18);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8879w(0) <= y_prenode_12_w(19);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8735w(0) <= y_prenode_12_w(1);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8887w(0) <= y_prenode_12_w(20);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8895w(0) <= y_prenode_12_w(21);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8903w(0) <= y_prenode_12_w(22);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8911w(0) <= y_prenode_12_w(23);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8919w(0) <= y_prenode_12_w(24);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8927w(0) <= y_prenode_12_w(25);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8935w(0) <= y_prenode_12_w(26);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8943w(0) <= y_prenode_12_w(27);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8951w(0) <= y_prenode_12_w(28);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8959w(0) <= y_prenode_12_w(29);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8743w(0) <= y_prenode_12_w(2);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8967w(0) <= y_prenode_12_w(30);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8975w(0) <= y_prenode_12_w(31);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8751w(0) <= y_prenode_12_w(3);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8759w(0) <= y_prenode_12_w(4);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8767w(0) <= y_prenode_12_w(5);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8775w(0) <= y_prenode_12_w(6);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8783w(0) <= y_prenode_12_w(7);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8791w(0) <= y_prenode_12_w(8);
	wire_ccc_cordic_m_w_y_prenode_12_w_range8799w(0) <= y_prenode_12_w(9);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9472w(0) <= y_prenode_13_w(0);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9553w(0) <= y_prenode_13_w(10);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9561w(0) <= y_prenode_13_w(11);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9569w(0) <= y_prenode_13_w(12);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9577w(0) <= y_prenode_13_w(13);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9585w(0) <= y_prenode_13_w(14);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9593w(0) <= y_prenode_13_w(15);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9601w(0) <= y_prenode_13_w(16);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9609w(0) <= y_prenode_13_w(17);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9617w(0) <= y_prenode_13_w(18);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9625w(0) <= y_prenode_13_w(19);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9481w(0) <= y_prenode_13_w(1);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9633w(0) <= y_prenode_13_w(20);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9641w(0) <= y_prenode_13_w(21);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9649w(0) <= y_prenode_13_w(22);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9657w(0) <= y_prenode_13_w(23);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9665w(0) <= y_prenode_13_w(24);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9673w(0) <= y_prenode_13_w(25);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9681w(0) <= y_prenode_13_w(26);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9689w(0) <= y_prenode_13_w(27);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9697w(0) <= y_prenode_13_w(28);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9705w(0) <= y_prenode_13_w(29);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9489w(0) <= y_prenode_13_w(2);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9713w(0) <= y_prenode_13_w(30);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9721w(0) <= y_prenode_13_w(31);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9497w(0) <= y_prenode_13_w(3);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9505w(0) <= y_prenode_13_w(4);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9513w(0) <= y_prenode_13_w(5);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9521w(0) <= y_prenode_13_w(6);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9529w(0) <= y_prenode_13_w(7);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9537w(0) <= y_prenode_13_w(8);
	wire_ccc_cordic_m_w_y_prenode_13_w_range9545w(0) <= y_prenode_13_w(9);
	wire_ccc_cordic_m_w_y_prenode_2_w_range991w(0) <= y_prenode_2_w(0);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1072w(0) <= y_prenode_2_w(10);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1080w(0) <= y_prenode_2_w(11);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1088w(0) <= y_prenode_2_w(12);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1096w(0) <= y_prenode_2_w(13);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1104w(0) <= y_prenode_2_w(14);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1112w(0) <= y_prenode_2_w(15);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1120w(0) <= y_prenode_2_w(16);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1128w(0) <= y_prenode_2_w(17);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1136w(0) <= y_prenode_2_w(18);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1144w(0) <= y_prenode_2_w(19);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1000w(0) <= y_prenode_2_w(1);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1152w(0) <= y_prenode_2_w(20);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1160w(0) <= y_prenode_2_w(21);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1168w(0) <= y_prenode_2_w(22);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1176w(0) <= y_prenode_2_w(23);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1184w(0) <= y_prenode_2_w(24);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1192w(0) <= y_prenode_2_w(25);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1200w(0) <= y_prenode_2_w(26);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1208w(0) <= y_prenode_2_w(27);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1216w(0) <= y_prenode_2_w(28);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1224w(0) <= y_prenode_2_w(29);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1008w(0) <= y_prenode_2_w(2);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1232w(0) <= y_prenode_2_w(30);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1240w(0) <= y_prenode_2_w(31);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1016w(0) <= y_prenode_2_w(3);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1024w(0) <= y_prenode_2_w(4);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1032w(0) <= y_prenode_2_w(5);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1040w(0) <= y_prenode_2_w(6);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1048w(0) <= y_prenode_2_w(7);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1056w(0) <= y_prenode_2_w(8);
	wire_ccc_cordic_m_w_y_prenode_2_w_range1064w(0) <= y_prenode_2_w(9);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1787w(0) <= y_prenode_3_w(0);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1868w(0) <= y_prenode_3_w(10);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1876w(0) <= y_prenode_3_w(11);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1884w(0) <= y_prenode_3_w(12);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1892w(0) <= y_prenode_3_w(13);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1900w(0) <= y_prenode_3_w(14);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1908w(0) <= y_prenode_3_w(15);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1916w(0) <= y_prenode_3_w(16);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1924w(0) <= y_prenode_3_w(17);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1932w(0) <= y_prenode_3_w(18);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1940w(0) <= y_prenode_3_w(19);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1796w(0) <= y_prenode_3_w(1);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1948w(0) <= y_prenode_3_w(20);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1956w(0) <= y_prenode_3_w(21);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1964w(0) <= y_prenode_3_w(22);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1972w(0) <= y_prenode_3_w(23);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1980w(0) <= y_prenode_3_w(24);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1988w(0) <= y_prenode_3_w(25);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1996w(0) <= y_prenode_3_w(26);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2004w(0) <= y_prenode_3_w(27);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2012w(0) <= y_prenode_3_w(28);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2020w(0) <= y_prenode_3_w(29);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1804w(0) <= y_prenode_3_w(2);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2028w(0) <= y_prenode_3_w(30);
	wire_ccc_cordic_m_w_y_prenode_3_w_range2036w(0) <= y_prenode_3_w(31);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1812w(0) <= y_prenode_3_w(3);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1820w(0) <= y_prenode_3_w(4);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1828w(0) <= y_prenode_3_w(5);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1836w(0) <= y_prenode_3_w(6);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1844w(0) <= y_prenode_3_w(7);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1852w(0) <= y_prenode_3_w(8);
	wire_ccc_cordic_m_w_y_prenode_3_w_range1860w(0) <= y_prenode_3_w(9);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2578w(0) <= y_prenode_4_w(0);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2659w(0) <= y_prenode_4_w(10);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2667w(0) <= y_prenode_4_w(11);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2675w(0) <= y_prenode_4_w(12);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2683w(0) <= y_prenode_4_w(13);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2691w(0) <= y_prenode_4_w(14);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2699w(0) <= y_prenode_4_w(15);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2707w(0) <= y_prenode_4_w(16);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2715w(0) <= y_prenode_4_w(17);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2723w(0) <= y_prenode_4_w(18);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2731w(0) <= y_prenode_4_w(19);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2587w(0) <= y_prenode_4_w(1);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2739w(0) <= y_prenode_4_w(20);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2747w(0) <= y_prenode_4_w(21);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2755w(0) <= y_prenode_4_w(22);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2763w(0) <= y_prenode_4_w(23);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2771w(0) <= y_prenode_4_w(24);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2779w(0) <= y_prenode_4_w(25);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2787w(0) <= y_prenode_4_w(26);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2795w(0) <= y_prenode_4_w(27);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2803w(0) <= y_prenode_4_w(28);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2811w(0) <= y_prenode_4_w(29);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2595w(0) <= y_prenode_4_w(2);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2819w(0) <= y_prenode_4_w(30);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2827w(0) <= y_prenode_4_w(31);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2603w(0) <= y_prenode_4_w(3);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2611w(0) <= y_prenode_4_w(4);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2619w(0) <= y_prenode_4_w(5);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2627w(0) <= y_prenode_4_w(6);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2635w(0) <= y_prenode_4_w(7);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2643w(0) <= y_prenode_4_w(8);
	wire_ccc_cordic_m_w_y_prenode_4_w_range2651w(0) <= y_prenode_4_w(9);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3364w(0) <= y_prenode_5_w(0);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3445w(0) <= y_prenode_5_w(10);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3453w(0) <= y_prenode_5_w(11);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3461w(0) <= y_prenode_5_w(12);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3469w(0) <= y_prenode_5_w(13);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3477w(0) <= y_prenode_5_w(14);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3485w(0) <= y_prenode_5_w(15);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3493w(0) <= y_prenode_5_w(16);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3501w(0) <= y_prenode_5_w(17);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3509w(0) <= y_prenode_5_w(18);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3517w(0) <= y_prenode_5_w(19);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3373w(0) <= y_prenode_5_w(1);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3525w(0) <= y_prenode_5_w(20);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3533w(0) <= y_prenode_5_w(21);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3541w(0) <= y_prenode_5_w(22);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3549w(0) <= y_prenode_5_w(23);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3557w(0) <= y_prenode_5_w(24);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3565w(0) <= y_prenode_5_w(25);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3573w(0) <= y_prenode_5_w(26);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3581w(0) <= y_prenode_5_w(27);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3589w(0) <= y_prenode_5_w(28);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3597w(0) <= y_prenode_5_w(29);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3381w(0) <= y_prenode_5_w(2);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3605w(0) <= y_prenode_5_w(30);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3613w(0) <= y_prenode_5_w(31);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3389w(0) <= y_prenode_5_w(3);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3397w(0) <= y_prenode_5_w(4);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3405w(0) <= y_prenode_5_w(5);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3413w(0) <= y_prenode_5_w(6);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3421w(0) <= y_prenode_5_w(7);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3429w(0) <= y_prenode_5_w(8);
	wire_ccc_cordic_m_w_y_prenode_5_w_range3437w(0) <= y_prenode_5_w(9);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4145w(0) <= y_prenode_6_w(0);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4226w(0) <= y_prenode_6_w(10);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4234w(0) <= y_prenode_6_w(11);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4242w(0) <= y_prenode_6_w(12);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4250w(0) <= y_prenode_6_w(13);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4258w(0) <= y_prenode_6_w(14);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4266w(0) <= y_prenode_6_w(15);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4274w(0) <= y_prenode_6_w(16);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4282w(0) <= y_prenode_6_w(17);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4290w(0) <= y_prenode_6_w(18);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4298w(0) <= y_prenode_6_w(19);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4154w(0) <= y_prenode_6_w(1);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4306w(0) <= y_prenode_6_w(20);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4314w(0) <= y_prenode_6_w(21);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4322w(0) <= y_prenode_6_w(22);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4330w(0) <= y_prenode_6_w(23);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4338w(0) <= y_prenode_6_w(24);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4346w(0) <= y_prenode_6_w(25);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4354w(0) <= y_prenode_6_w(26);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4362w(0) <= y_prenode_6_w(27);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4370w(0) <= y_prenode_6_w(28);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4378w(0) <= y_prenode_6_w(29);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4162w(0) <= y_prenode_6_w(2);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4386w(0) <= y_prenode_6_w(30);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4394w(0) <= y_prenode_6_w(31);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4170w(0) <= y_prenode_6_w(3);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4178w(0) <= y_prenode_6_w(4);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4186w(0) <= y_prenode_6_w(5);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4194w(0) <= y_prenode_6_w(6);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4202w(0) <= y_prenode_6_w(7);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4210w(0) <= y_prenode_6_w(8);
	wire_ccc_cordic_m_w_y_prenode_6_w_range4218w(0) <= y_prenode_6_w(9);
	wire_ccc_cordic_m_w_y_prenode_7_w_range4921w(0) <= y_prenode_7_w(0);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5002w(0) <= y_prenode_7_w(10);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5010w(0) <= y_prenode_7_w(11);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5018w(0) <= y_prenode_7_w(12);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5026w(0) <= y_prenode_7_w(13);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5034w(0) <= y_prenode_7_w(14);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5042w(0) <= y_prenode_7_w(15);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5050w(0) <= y_prenode_7_w(16);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5058w(0) <= y_prenode_7_w(17);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5066w(0) <= y_prenode_7_w(18);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5074w(0) <= y_prenode_7_w(19);
	wire_ccc_cordic_m_w_y_prenode_7_w_range4930w(0) <= y_prenode_7_w(1);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5082w(0) <= y_prenode_7_w(20);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5090w(0) <= y_prenode_7_w(21);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5098w(0) <= y_prenode_7_w(22);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5106w(0) <= y_prenode_7_w(23);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5114w(0) <= y_prenode_7_w(24);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5122w(0) <= y_prenode_7_w(25);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5130w(0) <= y_prenode_7_w(26);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5138w(0) <= y_prenode_7_w(27);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5146w(0) <= y_prenode_7_w(28);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5154w(0) <= y_prenode_7_w(29);
	wire_ccc_cordic_m_w_y_prenode_7_w_range4938w(0) <= y_prenode_7_w(2);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5162w(0) <= y_prenode_7_w(30);
	wire_ccc_cordic_m_w_y_prenode_7_w_range5170w(0) <= y_prenode_7_w(31);
	wire_ccc_cordic_m_w_y_prenode_7_w_range4946w(0) <= y_prenode_7_w(3);
	wire_ccc_cordic_m_w_y_prenode_7_w_range4954w(0) <= y_prenode_7_w(4);
	wire_ccc_cordic_m_w_y_prenode_7_w_range4962w(0) <= y_prenode_7_w(5);
	wire_ccc_cordic_m_w_y_prenode_7_w_range4970w(0) <= y_prenode_7_w(6);
	wire_ccc_cordic_m_w_y_prenode_7_w_range4978w(0) <= y_prenode_7_w(7);
	wire_ccc_cordic_m_w_y_prenode_7_w_range4986w(0) <= y_prenode_7_w(8);
	wire_ccc_cordic_m_w_y_prenode_7_w_range4994w(0) <= y_prenode_7_w(9);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5692w(0) <= y_prenode_8_w(0);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5773w(0) <= y_prenode_8_w(10);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5781w(0) <= y_prenode_8_w(11);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5789w(0) <= y_prenode_8_w(12);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5797w(0) <= y_prenode_8_w(13);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5805w(0) <= y_prenode_8_w(14);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5813w(0) <= y_prenode_8_w(15);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5821w(0) <= y_prenode_8_w(16);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5829w(0) <= y_prenode_8_w(17);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5837w(0) <= y_prenode_8_w(18);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5845w(0) <= y_prenode_8_w(19);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5701w(0) <= y_prenode_8_w(1);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5853w(0) <= y_prenode_8_w(20);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5861w(0) <= y_prenode_8_w(21);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5869w(0) <= y_prenode_8_w(22);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5877w(0) <= y_prenode_8_w(23);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5885w(0) <= y_prenode_8_w(24);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5893w(0) <= y_prenode_8_w(25);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5901w(0) <= y_prenode_8_w(26);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5909w(0) <= y_prenode_8_w(27);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5917w(0) <= y_prenode_8_w(28);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5925w(0) <= y_prenode_8_w(29);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5709w(0) <= y_prenode_8_w(2);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5933w(0) <= y_prenode_8_w(30);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5941w(0) <= y_prenode_8_w(31);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5717w(0) <= y_prenode_8_w(3);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5725w(0) <= y_prenode_8_w(4);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5733w(0) <= y_prenode_8_w(5);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5741w(0) <= y_prenode_8_w(6);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5749w(0) <= y_prenode_8_w(7);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5757w(0) <= y_prenode_8_w(8);
	wire_ccc_cordic_m_w_y_prenode_8_w_range5765w(0) <= y_prenode_8_w(9);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6458w(0) <= y_prenode_9_w(0);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6539w(0) <= y_prenode_9_w(10);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6547w(0) <= y_prenode_9_w(11);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6555w(0) <= y_prenode_9_w(12);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6563w(0) <= y_prenode_9_w(13);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6571w(0) <= y_prenode_9_w(14);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6579w(0) <= y_prenode_9_w(15);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6587w(0) <= y_prenode_9_w(16);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6595w(0) <= y_prenode_9_w(17);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6603w(0) <= y_prenode_9_w(18);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6611w(0) <= y_prenode_9_w(19);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6467w(0) <= y_prenode_9_w(1);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6619w(0) <= y_prenode_9_w(20);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6627w(0) <= y_prenode_9_w(21);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6635w(0) <= y_prenode_9_w(22);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6643w(0) <= y_prenode_9_w(23);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6651w(0) <= y_prenode_9_w(24);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6659w(0) <= y_prenode_9_w(25);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6667w(0) <= y_prenode_9_w(26);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6675w(0) <= y_prenode_9_w(27);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6683w(0) <= y_prenode_9_w(28);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6691w(0) <= y_prenode_9_w(29);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6475w(0) <= y_prenode_9_w(2);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6699w(0) <= y_prenode_9_w(30);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6707w(0) <= y_prenode_9_w(31);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6483w(0) <= y_prenode_9_w(3);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6491w(0) <= y_prenode_9_w(4);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6499w(0) <= y_prenode_9_w(5);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6507w(0) <= y_prenode_9_w(6);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6515w(0) <= y_prenode_9_w(7);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6523w(0) <= y_prenode_9_w(8);
	wire_ccc_cordic_m_w_y_prenode_9_w_range6531w(0) <= y_prenode_9_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7021w(0) <= y_prenodeone_10_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7080w(0) <= y_prenodeone_10_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7086w(0) <= y_prenodeone_10_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7092w(0) <= y_prenodeone_10_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7098w(0) <= y_prenodeone_10_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7104w(0) <= y_prenodeone_10_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7110w(0) <= y_prenodeone_10_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7116w(0) <= y_prenodeone_10_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7122w(0) <= y_prenodeone_10_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7128w(0) <= y_prenodeone_10_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7134w(0) <= y_prenodeone_10_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7026w(0) <= y_prenodeone_10_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7140w(0) <= y_prenodeone_10_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7146w(0) <= y_prenodeone_10_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7149w(0) <= y_prenodeone_10_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range6973w(0) <= y_prenodeone_10_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range6976w(0) <= y_prenodeone_10_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range6978w(0) <= y_prenodeone_10_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range6980w(0) <= y_prenodeone_10_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range6982w(0) <= y_prenodeone_10_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range6984w(0) <= y_prenodeone_10_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range6986w(0) <= y_prenodeone_10_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7032w(0) <= y_prenodeone_10_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range6988w(0) <= y_prenodeone_10_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range6990w(0) <= y_prenodeone_10_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7038w(0) <= y_prenodeone_10_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7044w(0) <= y_prenodeone_10_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7050w(0) <= y_prenodeone_10_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7056w(0) <= y_prenodeone_10_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7062w(0) <= y_prenodeone_10_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7068w(0) <= y_prenodeone_10_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_10_w_range7074w(0) <= y_prenodeone_10_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7786w(0) <= y_prenodeone_11_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7845w(0) <= y_prenodeone_11_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7851w(0) <= y_prenodeone_11_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7857w(0) <= y_prenodeone_11_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7863w(0) <= y_prenodeone_11_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7869w(0) <= y_prenodeone_11_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7875w(0) <= y_prenodeone_11_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7881w(0) <= y_prenodeone_11_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7887w(0) <= y_prenodeone_11_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7893w(0) <= y_prenodeone_11_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7899w(0) <= y_prenodeone_11_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7791w(0) <= y_prenodeone_11_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7905w(0) <= y_prenodeone_11_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7908w(0) <= y_prenodeone_11_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7734w(0) <= y_prenodeone_11_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7737w(0) <= y_prenodeone_11_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7739w(0) <= y_prenodeone_11_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7741w(0) <= y_prenodeone_11_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7743w(0) <= y_prenodeone_11_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7745w(0) <= y_prenodeone_11_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7747w(0) <= y_prenodeone_11_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7749w(0) <= y_prenodeone_11_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7797w(0) <= y_prenodeone_11_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7751w(0) <= y_prenodeone_11_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7753w(0) <= y_prenodeone_11_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7803w(0) <= y_prenodeone_11_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7809w(0) <= y_prenodeone_11_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7815w(0) <= y_prenodeone_11_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7821w(0) <= y_prenodeone_11_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7827w(0) <= y_prenodeone_11_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7833w(0) <= y_prenodeone_11_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_11_w_range7839w(0) <= y_prenodeone_11_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8546w(0) <= y_prenodeone_12_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8605w(0) <= y_prenodeone_12_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8611w(0) <= y_prenodeone_12_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8617w(0) <= y_prenodeone_12_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8623w(0) <= y_prenodeone_12_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8629w(0) <= y_prenodeone_12_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8635w(0) <= y_prenodeone_12_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8641w(0) <= y_prenodeone_12_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8647w(0) <= y_prenodeone_12_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8653w(0) <= y_prenodeone_12_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8659w(0) <= y_prenodeone_12_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8551w(0) <= y_prenodeone_12_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8662w(0) <= y_prenodeone_12_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8490w(0) <= y_prenodeone_12_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8493w(0) <= y_prenodeone_12_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8495w(0) <= y_prenodeone_12_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8497w(0) <= y_prenodeone_12_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8499w(0) <= y_prenodeone_12_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8501w(0) <= y_prenodeone_12_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8503w(0) <= y_prenodeone_12_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8505w(0) <= y_prenodeone_12_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8507w(0) <= y_prenodeone_12_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8557w(0) <= y_prenodeone_12_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8509w(0) <= y_prenodeone_12_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8511w(0) <= y_prenodeone_12_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8563w(0) <= y_prenodeone_12_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8569w(0) <= y_prenodeone_12_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8575w(0) <= y_prenodeone_12_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8581w(0) <= y_prenodeone_12_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8587w(0) <= y_prenodeone_12_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8593w(0) <= y_prenodeone_12_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_12_w_range8599w(0) <= y_prenodeone_12_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9301w(0) <= y_prenodeone_13_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9360w(0) <= y_prenodeone_13_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9366w(0) <= y_prenodeone_13_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9372w(0) <= y_prenodeone_13_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9378w(0) <= y_prenodeone_13_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9384w(0) <= y_prenodeone_13_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9390w(0) <= y_prenodeone_13_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9396w(0) <= y_prenodeone_13_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9402w(0) <= y_prenodeone_13_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9408w(0) <= y_prenodeone_13_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9411w(0) <= y_prenodeone_13_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9306w(0) <= y_prenodeone_13_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9241w(0) <= y_prenodeone_13_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9244w(0) <= y_prenodeone_13_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9246w(0) <= y_prenodeone_13_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9248w(0) <= y_prenodeone_13_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9250w(0) <= y_prenodeone_13_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9252w(0) <= y_prenodeone_13_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9254w(0) <= y_prenodeone_13_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9256w(0) <= y_prenodeone_13_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9258w(0) <= y_prenodeone_13_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9260w(0) <= y_prenodeone_13_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9312w(0) <= y_prenodeone_13_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9262w(0) <= y_prenodeone_13_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9264w(0) <= y_prenodeone_13_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9318w(0) <= y_prenodeone_13_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9324w(0) <= y_prenodeone_13_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9330w(0) <= y_prenodeone_13_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9336w(0) <= y_prenodeone_13_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9342w(0) <= y_prenodeone_13_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9348w(0) <= y_prenodeone_13_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_13_w_range9354w(0) <= y_prenodeone_13_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range721w(0) <= y_prenodeone_2_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range780w(0) <= y_prenodeone_2_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range786w(0) <= y_prenodeone_2_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range792w(0) <= y_prenodeone_2_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range798w(0) <= y_prenodeone_2_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range804w(0) <= y_prenodeone_2_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range810w(0) <= y_prenodeone_2_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range816w(0) <= y_prenodeone_2_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range822w(0) <= y_prenodeone_2_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range828w(0) <= y_prenodeone_2_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range834w(0) <= y_prenodeone_2_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range726w(0) <= y_prenodeone_2_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range840w(0) <= y_prenodeone_2_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range846w(0) <= y_prenodeone_2_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range852w(0) <= y_prenodeone_2_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range858w(0) <= y_prenodeone_2_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range864w(0) <= y_prenodeone_2_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range870w(0) <= y_prenodeone_2_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range876w(0) <= y_prenodeone_2_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range882w(0) <= y_prenodeone_2_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range888w(0) <= y_prenodeone_2_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range894w(0) <= y_prenodeone_2_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range732w(0) <= y_prenodeone_2_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range897w(0) <= y_prenodeone_2_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range705w(0) <= y_prenodeone_2_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range738w(0) <= y_prenodeone_2_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range744w(0) <= y_prenodeone_2_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range750w(0) <= y_prenodeone_2_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range756w(0) <= y_prenodeone_2_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range762w(0) <= y_prenodeone_2_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range768w(0) <= y_prenodeone_2_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_2_w_range774w(0) <= y_prenodeone_2_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1526w(0) <= y_prenodeone_3_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1585w(0) <= y_prenodeone_3_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1591w(0) <= y_prenodeone_3_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1597w(0) <= y_prenodeone_3_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1603w(0) <= y_prenodeone_3_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1609w(0) <= y_prenodeone_3_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1615w(0) <= y_prenodeone_3_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1621w(0) <= y_prenodeone_3_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1627w(0) <= y_prenodeone_3_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1633w(0) <= y_prenodeone_3_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1639w(0) <= y_prenodeone_3_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1531w(0) <= y_prenodeone_3_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1645w(0) <= y_prenodeone_3_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1651w(0) <= y_prenodeone_3_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1657w(0) <= y_prenodeone_3_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1663w(0) <= y_prenodeone_3_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1669w(0) <= y_prenodeone_3_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1675w(0) <= y_prenodeone_3_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1681w(0) <= y_prenodeone_3_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1687w(0) <= y_prenodeone_3_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1693w(0) <= y_prenodeone_3_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1696w(0) <= y_prenodeone_3_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1537w(0) <= y_prenodeone_3_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1506w(0) <= y_prenodeone_3_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1509w(0) <= y_prenodeone_3_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1543w(0) <= y_prenodeone_3_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1549w(0) <= y_prenodeone_3_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1555w(0) <= y_prenodeone_3_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1561w(0) <= y_prenodeone_3_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1567w(0) <= y_prenodeone_3_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1573w(0) <= y_prenodeone_3_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_3_w_range1579w(0) <= y_prenodeone_3_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2326w(0) <= y_prenodeone_4_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2385w(0) <= y_prenodeone_4_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2391w(0) <= y_prenodeone_4_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2397w(0) <= y_prenodeone_4_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2403w(0) <= y_prenodeone_4_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2409w(0) <= y_prenodeone_4_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2415w(0) <= y_prenodeone_4_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2421w(0) <= y_prenodeone_4_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2427w(0) <= y_prenodeone_4_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2433w(0) <= y_prenodeone_4_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2439w(0) <= y_prenodeone_4_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2331w(0) <= y_prenodeone_4_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2445w(0) <= y_prenodeone_4_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2451w(0) <= y_prenodeone_4_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2457w(0) <= y_prenodeone_4_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2463w(0) <= y_prenodeone_4_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2469w(0) <= y_prenodeone_4_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2475w(0) <= y_prenodeone_4_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2481w(0) <= y_prenodeone_4_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2487w(0) <= y_prenodeone_4_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2490w(0) <= y_prenodeone_4_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2302w(0) <= y_prenodeone_4_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2337w(0) <= y_prenodeone_4_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2305w(0) <= y_prenodeone_4_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2307w(0) <= y_prenodeone_4_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2343w(0) <= y_prenodeone_4_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2349w(0) <= y_prenodeone_4_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2355w(0) <= y_prenodeone_4_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2361w(0) <= y_prenodeone_4_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2367w(0) <= y_prenodeone_4_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2373w(0) <= y_prenodeone_4_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_4_w_range2379w(0) <= y_prenodeone_4_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3121w(0) <= y_prenodeone_5_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3180w(0) <= y_prenodeone_5_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3186w(0) <= y_prenodeone_5_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3192w(0) <= y_prenodeone_5_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3198w(0) <= y_prenodeone_5_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3204w(0) <= y_prenodeone_5_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3210w(0) <= y_prenodeone_5_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3216w(0) <= y_prenodeone_5_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3222w(0) <= y_prenodeone_5_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3228w(0) <= y_prenodeone_5_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3234w(0) <= y_prenodeone_5_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3126w(0) <= y_prenodeone_5_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3240w(0) <= y_prenodeone_5_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3246w(0) <= y_prenodeone_5_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3252w(0) <= y_prenodeone_5_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3258w(0) <= y_prenodeone_5_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3264w(0) <= y_prenodeone_5_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3270w(0) <= y_prenodeone_5_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3276w(0) <= y_prenodeone_5_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3279w(0) <= y_prenodeone_5_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3093w(0) <= y_prenodeone_5_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3096w(0) <= y_prenodeone_5_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3132w(0) <= y_prenodeone_5_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3098w(0) <= y_prenodeone_5_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3100w(0) <= y_prenodeone_5_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3138w(0) <= y_prenodeone_5_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3144w(0) <= y_prenodeone_5_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3150w(0) <= y_prenodeone_5_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3156w(0) <= y_prenodeone_5_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3162w(0) <= y_prenodeone_5_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3168w(0) <= y_prenodeone_5_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_5_w_range3174w(0) <= y_prenodeone_5_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3911w(0) <= y_prenodeone_6_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3970w(0) <= y_prenodeone_6_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3976w(0) <= y_prenodeone_6_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3982w(0) <= y_prenodeone_6_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3988w(0) <= y_prenodeone_6_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3994w(0) <= y_prenodeone_6_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4000w(0) <= y_prenodeone_6_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4006w(0) <= y_prenodeone_6_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4012w(0) <= y_prenodeone_6_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4018w(0) <= y_prenodeone_6_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4024w(0) <= y_prenodeone_6_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3916w(0) <= y_prenodeone_6_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4030w(0) <= y_prenodeone_6_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4036w(0) <= y_prenodeone_6_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4042w(0) <= y_prenodeone_6_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4048w(0) <= y_prenodeone_6_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4054w(0) <= y_prenodeone_6_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4060w(0) <= y_prenodeone_6_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range4063w(0) <= y_prenodeone_6_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3879w(0) <= y_prenodeone_6_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3882w(0) <= y_prenodeone_6_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3884w(0) <= y_prenodeone_6_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3922w(0) <= y_prenodeone_6_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3886w(0) <= y_prenodeone_6_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3888w(0) <= y_prenodeone_6_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3928w(0) <= y_prenodeone_6_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3934w(0) <= y_prenodeone_6_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3940w(0) <= y_prenodeone_6_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3946w(0) <= y_prenodeone_6_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3952w(0) <= y_prenodeone_6_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3958w(0) <= y_prenodeone_6_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_6_w_range3964w(0) <= y_prenodeone_6_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4696w(0) <= y_prenodeone_7_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4755w(0) <= y_prenodeone_7_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4761w(0) <= y_prenodeone_7_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4767w(0) <= y_prenodeone_7_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4773w(0) <= y_prenodeone_7_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4779w(0) <= y_prenodeone_7_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4785w(0) <= y_prenodeone_7_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4791w(0) <= y_prenodeone_7_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4797w(0) <= y_prenodeone_7_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4803w(0) <= y_prenodeone_7_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4809w(0) <= y_prenodeone_7_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4701w(0) <= y_prenodeone_7_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4815w(0) <= y_prenodeone_7_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4821w(0) <= y_prenodeone_7_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4827w(0) <= y_prenodeone_7_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4833w(0) <= y_prenodeone_7_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4839w(0) <= y_prenodeone_7_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4842w(0) <= y_prenodeone_7_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4660w(0) <= y_prenodeone_7_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4663w(0) <= y_prenodeone_7_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4665w(0) <= y_prenodeone_7_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4667w(0) <= y_prenodeone_7_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4707w(0) <= y_prenodeone_7_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4669w(0) <= y_prenodeone_7_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4671w(0) <= y_prenodeone_7_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4713w(0) <= y_prenodeone_7_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4719w(0) <= y_prenodeone_7_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4725w(0) <= y_prenodeone_7_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4731w(0) <= y_prenodeone_7_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4737w(0) <= y_prenodeone_7_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4743w(0) <= y_prenodeone_7_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_7_w_range4749w(0) <= y_prenodeone_7_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5476w(0) <= y_prenodeone_8_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5535w(0) <= y_prenodeone_8_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5541w(0) <= y_prenodeone_8_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5547w(0) <= y_prenodeone_8_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5553w(0) <= y_prenodeone_8_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5559w(0) <= y_prenodeone_8_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5565w(0) <= y_prenodeone_8_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5571w(0) <= y_prenodeone_8_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5577w(0) <= y_prenodeone_8_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5583w(0) <= y_prenodeone_8_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5589w(0) <= y_prenodeone_8_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5481w(0) <= y_prenodeone_8_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5595w(0) <= y_prenodeone_8_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5601w(0) <= y_prenodeone_8_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5607w(0) <= y_prenodeone_8_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5613w(0) <= y_prenodeone_8_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5616w(0) <= y_prenodeone_8_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5436w(0) <= y_prenodeone_8_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5439w(0) <= y_prenodeone_8_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5441w(0) <= y_prenodeone_8_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5443w(0) <= y_prenodeone_8_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5445w(0) <= y_prenodeone_8_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5487w(0) <= y_prenodeone_8_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5447w(0) <= y_prenodeone_8_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5449w(0) <= y_prenodeone_8_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5493w(0) <= y_prenodeone_8_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5499w(0) <= y_prenodeone_8_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5505w(0) <= y_prenodeone_8_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5511w(0) <= y_prenodeone_8_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5517w(0) <= y_prenodeone_8_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5523w(0) <= y_prenodeone_8_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_8_w_range5529w(0) <= y_prenodeone_8_w(9);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6251w(0) <= y_prenodeone_9_w(0);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6310w(0) <= y_prenodeone_9_w(10);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6316w(0) <= y_prenodeone_9_w(11);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6322w(0) <= y_prenodeone_9_w(12);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6328w(0) <= y_prenodeone_9_w(13);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6334w(0) <= y_prenodeone_9_w(14);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6340w(0) <= y_prenodeone_9_w(15);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6346w(0) <= y_prenodeone_9_w(16);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6352w(0) <= y_prenodeone_9_w(17);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6358w(0) <= y_prenodeone_9_w(18);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6364w(0) <= y_prenodeone_9_w(19);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6256w(0) <= y_prenodeone_9_w(1);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6370w(0) <= y_prenodeone_9_w(20);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6376w(0) <= y_prenodeone_9_w(21);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6382w(0) <= y_prenodeone_9_w(22);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6385w(0) <= y_prenodeone_9_w(23);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6207w(0) <= y_prenodeone_9_w(24);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6210w(0) <= y_prenodeone_9_w(25);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6212w(0) <= y_prenodeone_9_w(26);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6214w(0) <= y_prenodeone_9_w(27);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6216w(0) <= y_prenodeone_9_w(28);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6218w(0) <= y_prenodeone_9_w(29);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6262w(0) <= y_prenodeone_9_w(2);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6220w(0) <= y_prenodeone_9_w(30);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6222w(0) <= y_prenodeone_9_w(31);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6268w(0) <= y_prenodeone_9_w(3);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6274w(0) <= y_prenodeone_9_w(4);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6280w(0) <= y_prenodeone_9_w(5);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6286w(0) <= y_prenodeone_9_w(6);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6292w(0) <= y_prenodeone_9_w(7);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6298w(0) <= y_prenodeone_9_w(8);
	wire_ccc_cordic_m_w_y_prenodeone_9_w_range6304w(0) <= y_prenodeone_9_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7152w(0) <= y_prenodetwo_10_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7181w(0) <= y_prenodetwo_10_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7184w(0) <= y_prenodetwo_10_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7187w(0) <= y_prenodetwo_10_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7190w(0) <= y_prenodetwo_10_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7193w(0) <= y_prenodetwo_10_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7196w(0) <= y_prenodetwo_10_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7199w(0) <= y_prenodetwo_10_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7202w(0) <= y_prenodetwo_10_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7205w(0) <= y_prenodetwo_10_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7208w(0) <= y_prenodetwo_10_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7154w(0) <= y_prenodetwo_10_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range6993w(0) <= y_prenodetwo_10_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range6996w(0) <= y_prenodetwo_10_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range6998w(0) <= y_prenodetwo_10_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7000w(0) <= y_prenodetwo_10_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7002w(0) <= y_prenodetwo_10_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7004w(0) <= y_prenodetwo_10_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7006w(0) <= y_prenodetwo_10_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7008w(0) <= y_prenodetwo_10_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7010w(0) <= y_prenodetwo_10_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7012w(0) <= y_prenodetwo_10_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7157w(0) <= y_prenodetwo_10_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7014w(0) <= y_prenodetwo_10_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7016w(0) <= y_prenodetwo_10_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7160w(0) <= y_prenodetwo_10_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7163w(0) <= y_prenodetwo_10_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7166w(0) <= y_prenodetwo_10_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7169w(0) <= y_prenodetwo_10_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7172w(0) <= y_prenodetwo_10_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7175w(0) <= y_prenodetwo_10_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_10_w_range7178w(0) <= y_prenodetwo_10_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7911w(0) <= y_prenodetwo_11_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7940w(0) <= y_prenodetwo_11_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7943w(0) <= y_prenodetwo_11_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7946w(0) <= y_prenodetwo_11_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7949w(0) <= y_prenodetwo_11_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7952w(0) <= y_prenodetwo_11_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7955w(0) <= y_prenodetwo_11_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7958w(0) <= y_prenodetwo_11_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7961w(0) <= y_prenodetwo_11_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7964w(0) <= y_prenodetwo_11_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7756w(0) <= y_prenodetwo_11_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7913w(0) <= y_prenodetwo_11_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7759w(0) <= y_prenodetwo_11_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7761w(0) <= y_prenodetwo_11_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7763w(0) <= y_prenodetwo_11_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7765w(0) <= y_prenodetwo_11_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7767w(0) <= y_prenodetwo_11_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7769w(0) <= y_prenodetwo_11_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7771w(0) <= y_prenodetwo_11_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7773w(0) <= y_prenodetwo_11_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7775w(0) <= y_prenodetwo_11_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7777w(0) <= y_prenodetwo_11_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7916w(0) <= y_prenodetwo_11_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7779w(0) <= y_prenodetwo_11_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7781w(0) <= y_prenodetwo_11_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7919w(0) <= y_prenodetwo_11_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7922w(0) <= y_prenodetwo_11_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7925w(0) <= y_prenodetwo_11_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7928w(0) <= y_prenodetwo_11_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7931w(0) <= y_prenodetwo_11_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7934w(0) <= y_prenodetwo_11_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_11_w_range7937w(0) <= y_prenodetwo_11_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8665w(0) <= y_prenodetwo_12_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8694w(0) <= y_prenodetwo_12_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8697w(0) <= y_prenodetwo_12_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8700w(0) <= y_prenodetwo_12_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8703w(0) <= y_prenodetwo_12_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8706w(0) <= y_prenodetwo_12_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8709w(0) <= y_prenodetwo_12_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8712w(0) <= y_prenodetwo_12_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8715w(0) <= y_prenodetwo_12_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8514w(0) <= y_prenodetwo_12_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8517w(0) <= y_prenodetwo_12_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8667w(0) <= y_prenodetwo_12_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8519w(0) <= y_prenodetwo_12_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8521w(0) <= y_prenodetwo_12_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8523w(0) <= y_prenodetwo_12_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8525w(0) <= y_prenodetwo_12_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8527w(0) <= y_prenodetwo_12_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8529w(0) <= y_prenodetwo_12_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8531w(0) <= y_prenodetwo_12_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8533w(0) <= y_prenodetwo_12_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8535w(0) <= y_prenodetwo_12_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8537w(0) <= y_prenodetwo_12_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8670w(0) <= y_prenodetwo_12_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8539w(0) <= y_prenodetwo_12_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8541w(0) <= y_prenodetwo_12_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8673w(0) <= y_prenodetwo_12_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8676w(0) <= y_prenodetwo_12_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8679w(0) <= y_prenodetwo_12_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8682w(0) <= y_prenodetwo_12_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8685w(0) <= y_prenodetwo_12_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8688w(0) <= y_prenodetwo_12_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_12_w_range8691w(0) <= y_prenodetwo_12_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9414w(0) <= y_prenodetwo_13_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9443w(0) <= y_prenodetwo_13_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9446w(0) <= y_prenodetwo_13_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9449w(0) <= y_prenodetwo_13_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9452w(0) <= y_prenodetwo_13_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9455w(0) <= y_prenodetwo_13_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9458w(0) <= y_prenodetwo_13_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9461w(0) <= y_prenodetwo_13_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9267w(0) <= y_prenodetwo_13_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9270w(0) <= y_prenodetwo_13_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9272w(0) <= y_prenodetwo_13_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9416w(0) <= y_prenodetwo_13_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9274w(0) <= y_prenodetwo_13_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9276w(0) <= y_prenodetwo_13_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9278w(0) <= y_prenodetwo_13_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9280w(0) <= y_prenodetwo_13_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9282w(0) <= y_prenodetwo_13_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9284w(0) <= y_prenodetwo_13_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9286w(0) <= y_prenodetwo_13_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9288w(0) <= y_prenodetwo_13_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9290w(0) <= y_prenodetwo_13_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9292w(0) <= y_prenodetwo_13_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9419w(0) <= y_prenodetwo_13_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9294w(0) <= y_prenodetwo_13_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9296w(0) <= y_prenodetwo_13_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9422w(0) <= y_prenodetwo_13_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9425w(0) <= y_prenodetwo_13_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9428w(0) <= y_prenodetwo_13_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9431w(0) <= y_prenodetwo_13_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9434w(0) <= y_prenodetwo_13_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9437w(0) <= y_prenodetwo_13_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_13_w_range9440w(0) <= y_prenodetwo_13_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range900w(0) <= y_prenodetwo_2_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range929w(0) <= y_prenodetwo_2_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range932w(0) <= y_prenodetwo_2_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range935w(0) <= y_prenodetwo_2_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range938w(0) <= y_prenodetwo_2_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range941w(0) <= y_prenodetwo_2_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range944w(0) <= y_prenodetwo_2_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range947w(0) <= y_prenodetwo_2_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range950w(0) <= y_prenodetwo_2_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range953w(0) <= y_prenodetwo_2_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range956w(0) <= y_prenodetwo_2_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range902w(0) <= y_prenodetwo_2_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range959w(0) <= y_prenodetwo_2_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range962w(0) <= y_prenodetwo_2_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range965w(0) <= y_prenodetwo_2_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range968w(0) <= y_prenodetwo_2_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range971w(0) <= y_prenodetwo_2_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range974w(0) <= y_prenodetwo_2_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range977w(0) <= y_prenodetwo_2_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range980w(0) <= y_prenodetwo_2_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range709w(0) <= y_prenodetwo_2_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range712w(0) <= y_prenodetwo_2_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range905w(0) <= y_prenodetwo_2_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range714w(0) <= y_prenodetwo_2_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range716w(0) <= y_prenodetwo_2_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range908w(0) <= y_prenodetwo_2_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range911w(0) <= y_prenodetwo_2_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range914w(0) <= y_prenodetwo_2_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range917w(0) <= y_prenodetwo_2_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range920w(0) <= y_prenodetwo_2_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range923w(0) <= y_prenodetwo_2_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_2_w_range926w(0) <= y_prenodetwo_2_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1699w(0) <= y_prenodetwo_3_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1728w(0) <= y_prenodetwo_3_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1731w(0) <= y_prenodetwo_3_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1734w(0) <= y_prenodetwo_3_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1737w(0) <= y_prenodetwo_3_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1740w(0) <= y_prenodetwo_3_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1743w(0) <= y_prenodetwo_3_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1746w(0) <= y_prenodetwo_3_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1749w(0) <= y_prenodetwo_3_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1752w(0) <= y_prenodetwo_3_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1755w(0) <= y_prenodetwo_3_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1701w(0) <= y_prenodetwo_3_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1758w(0) <= y_prenodetwo_3_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1761w(0) <= y_prenodetwo_3_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1764w(0) <= y_prenodetwo_3_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1767w(0) <= y_prenodetwo_3_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1770w(0) <= y_prenodetwo_3_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1773w(0) <= y_prenodetwo_3_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1776w(0) <= y_prenodetwo_3_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1512w(0) <= y_prenodetwo_3_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1515w(0) <= y_prenodetwo_3_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1517w(0) <= y_prenodetwo_3_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1704w(0) <= y_prenodetwo_3_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1519w(0) <= y_prenodetwo_3_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1521w(0) <= y_prenodetwo_3_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1707w(0) <= y_prenodetwo_3_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1710w(0) <= y_prenodetwo_3_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1713w(0) <= y_prenodetwo_3_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1716w(0) <= y_prenodetwo_3_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1719w(0) <= y_prenodetwo_3_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1722w(0) <= y_prenodetwo_3_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_3_w_range1725w(0) <= y_prenodetwo_3_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2493w(0) <= y_prenodetwo_4_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2522w(0) <= y_prenodetwo_4_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2525w(0) <= y_prenodetwo_4_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2528w(0) <= y_prenodetwo_4_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2531w(0) <= y_prenodetwo_4_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2534w(0) <= y_prenodetwo_4_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2537w(0) <= y_prenodetwo_4_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2540w(0) <= y_prenodetwo_4_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2543w(0) <= y_prenodetwo_4_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2546w(0) <= y_prenodetwo_4_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2549w(0) <= y_prenodetwo_4_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2495w(0) <= y_prenodetwo_4_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2552w(0) <= y_prenodetwo_4_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2555w(0) <= y_prenodetwo_4_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2558w(0) <= y_prenodetwo_4_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2561w(0) <= y_prenodetwo_4_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2564w(0) <= y_prenodetwo_4_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2567w(0) <= y_prenodetwo_4_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2310w(0) <= y_prenodetwo_4_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2313w(0) <= y_prenodetwo_4_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2315w(0) <= y_prenodetwo_4_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2317w(0) <= y_prenodetwo_4_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2498w(0) <= y_prenodetwo_4_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2319w(0) <= y_prenodetwo_4_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2321w(0) <= y_prenodetwo_4_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2501w(0) <= y_prenodetwo_4_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2504w(0) <= y_prenodetwo_4_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2507w(0) <= y_prenodetwo_4_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2510w(0) <= y_prenodetwo_4_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2513w(0) <= y_prenodetwo_4_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2516w(0) <= y_prenodetwo_4_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_4_w_range2519w(0) <= y_prenodetwo_4_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3282w(0) <= y_prenodetwo_5_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3311w(0) <= y_prenodetwo_5_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3314w(0) <= y_prenodetwo_5_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3317w(0) <= y_prenodetwo_5_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3320w(0) <= y_prenodetwo_5_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3323w(0) <= y_prenodetwo_5_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3326w(0) <= y_prenodetwo_5_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3329w(0) <= y_prenodetwo_5_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3332w(0) <= y_prenodetwo_5_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3335w(0) <= y_prenodetwo_5_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3338w(0) <= y_prenodetwo_5_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3284w(0) <= y_prenodetwo_5_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3341w(0) <= y_prenodetwo_5_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3344w(0) <= y_prenodetwo_5_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3347w(0) <= y_prenodetwo_5_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3350w(0) <= y_prenodetwo_5_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3353w(0) <= y_prenodetwo_5_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3103w(0) <= y_prenodetwo_5_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3106w(0) <= y_prenodetwo_5_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3108w(0) <= y_prenodetwo_5_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3110w(0) <= y_prenodetwo_5_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3112w(0) <= y_prenodetwo_5_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3287w(0) <= y_prenodetwo_5_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3114w(0) <= y_prenodetwo_5_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3116w(0) <= y_prenodetwo_5_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3290w(0) <= y_prenodetwo_5_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3293w(0) <= y_prenodetwo_5_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3296w(0) <= y_prenodetwo_5_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3299w(0) <= y_prenodetwo_5_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3302w(0) <= y_prenodetwo_5_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3305w(0) <= y_prenodetwo_5_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_5_w_range3308w(0) <= y_prenodetwo_5_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4066w(0) <= y_prenodetwo_6_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4095w(0) <= y_prenodetwo_6_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4098w(0) <= y_prenodetwo_6_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4101w(0) <= y_prenodetwo_6_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4104w(0) <= y_prenodetwo_6_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4107w(0) <= y_prenodetwo_6_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4110w(0) <= y_prenodetwo_6_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4113w(0) <= y_prenodetwo_6_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4116w(0) <= y_prenodetwo_6_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4119w(0) <= y_prenodetwo_6_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4122w(0) <= y_prenodetwo_6_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4068w(0) <= y_prenodetwo_6_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4125w(0) <= y_prenodetwo_6_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4128w(0) <= y_prenodetwo_6_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4131w(0) <= y_prenodetwo_6_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4134w(0) <= y_prenodetwo_6_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3891w(0) <= y_prenodetwo_6_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3894w(0) <= y_prenodetwo_6_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3896w(0) <= y_prenodetwo_6_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3898w(0) <= y_prenodetwo_6_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3900w(0) <= y_prenodetwo_6_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3902w(0) <= y_prenodetwo_6_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4071w(0) <= y_prenodetwo_6_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3904w(0) <= y_prenodetwo_6_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range3906w(0) <= y_prenodetwo_6_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4074w(0) <= y_prenodetwo_6_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4077w(0) <= y_prenodetwo_6_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4080w(0) <= y_prenodetwo_6_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4083w(0) <= y_prenodetwo_6_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4086w(0) <= y_prenodetwo_6_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4089w(0) <= y_prenodetwo_6_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_6_w_range4092w(0) <= y_prenodetwo_6_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4845w(0) <= y_prenodetwo_7_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4874w(0) <= y_prenodetwo_7_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4877w(0) <= y_prenodetwo_7_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4880w(0) <= y_prenodetwo_7_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4883w(0) <= y_prenodetwo_7_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4886w(0) <= y_prenodetwo_7_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4889w(0) <= y_prenodetwo_7_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4892w(0) <= y_prenodetwo_7_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4895w(0) <= y_prenodetwo_7_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4898w(0) <= y_prenodetwo_7_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4901w(0) <= y_prenodetwo_7_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4847w(0) <= y_prenodetwo_7_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4904w(0) <= y_prenodetwo_7_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4907w(0) <= y_prenodetwo_7_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4910w(0) <= y_prenodetwo_7_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4674w(0) <= y_prenodetwo_7_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4677w(0) <= y_prenodetwo_7_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4679w(0) <= y_prenodetwo_7_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4681w(0) <= y_prenodetwo_7_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4683w(0) <= y_prenodetwo_7_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4685w(0) <= y_prenodetwo_7_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4687w(0) <= y_prenodetwo_7_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4850w(0) <= y_prenodetwo_7_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4689w(0) <= y_prenodetwo_7_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4691w(0) <= y_prenodetwo_7_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4853w(0) <= y_prenodetwo_7_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4856w(0) <= y_prenodetwo_7_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4859w(0) <= y_prenodetwo_7_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4862w(0) <= y_prenodetwo_7_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4865w(0) <= y_prenodetwo_7_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4868w(0) <= y_prenodetwo_7_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_7_w_range4871w(0) <= y_prenodetwo_7_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5619w(0) <= y_prenodetwo_8_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5648w(0) <= y_prenodetwo_8_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5651w(0) <= y_prenodetwo_8_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5654w(0) <= y_prenodetwo_8_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5657w(0) <= y_prenodetwo_8_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5660w(0) <= y_prenodetwo_8_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5663w(0) <= y_prenodetwo_8_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5666w(0) <= y_prenodetwo_8_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5669w(0) <= y_prenodetwo_8_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5672w(0) <= y_prenodetwo_8_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5675w(0) <= y_prenodetwo_8_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5621w(0) <= y_prenodetwo_8_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5678w(0) <= y_prenodetwo_8_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5681w(0) <= y_prenodetwo_8_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5452w(0) <= y_prenodetwo_8_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5455w(0) <= y_prenodetwo_8_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5457w(0) <= y_prenodetwo_8_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5459w(0) <= y_prenodetwo_8_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5461w(0) <= y_prenodetwo_8_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5463w(0) <= y_prenodetwo_8_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5465w(0) <= y_prenodetwo_8_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5467w(0) <= y_prenodetwo_8_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5624w(0) <= y_prenodetwo_8_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5469w(0) <= y_prenodetwo_8_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5471w(0) <= y_prenodetwo_8_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5627w(0) <= y_prenodetwo_8_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5630w(0) <= y_prenodetwo_8_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5633w(0) <= y_prenodetwo_8_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5636w(0) <= y_prenodetwo_8_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5639w(0) <= y_prenodetwo_8_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5642w(0) <= y_prenodetwo_8_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_8_w_range5645w(0) <= y_prenodetwo_8_w(9);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6388w(0) <= y_prenodetwo_9_w(0);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6417w(0) <= y_prenodetwo_9_w(10);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6420w(0) <= y_prenodetwo_9_w(11);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6423w(0) <= y_prenodetwo_9_w(12);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6426w(0) <= y_prenodetwo_9_w(13);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6429w(0) <= y_prenodetwo_9_w(14);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6432w(0) <= y_prenodetwo_9_w(15);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6435w(0) <= y_prenodetwo_9_w(16);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6438w(0) <= y_prenodetwo_9_w(17);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6441w(0) <= y_prenodetwo_9_w(18);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6444w(0) <= y_prenodetwo_9_w(19);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6390w(0) <= y_prenodetwo_9_w(1);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6447w(0) <= y_prenodetwo_9_w(20);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6225w(0) <= y_prenodetwo_9_w(21);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6228w(0) <= y_prenodetwo_9_w(22);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6230w(0) <= y_prenodetwo_9_w(23);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6232w(0) <= y_prenodetwo_9_w(24);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6234w(0) <= y_prenodetwo_9_w(25);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6236w(0) <= y_prenodetwo_9_w(26);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6238w(0) <= y_prenodetwo_9_w(27);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6240w(0) <= y_prenodetwo_9_w(28);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6242w(0) <= y_prenodetwo_9_w(29);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6393w(0) <= y_prenodetwo_9_w(2);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6244w(0) <= y_prenodetwo_9_w(30);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6246w(0) <= y_prenodetwo_9_w(31);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6396w(0) <= y_prenodetwo_9_w(3);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6399w(0) <= y_prenodetwo_9_w(4);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6402w(0) <= y_prenodetwo_9_w(5);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6405w(0) <= y_prenodetwo_9_w(6);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6408w(0) <= y_prenodetwo_9_w(7);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6411w(0) <= y_prenodetwo_9_w(8);
	wire_ccc_cordic_m_w_y_prenodetwo_9_w_range6414w(0) <= y_prenodetwo_9_w(9);
	cata_0_cordic_atan :  coshw_altfp_sincos_cordic_atan_35b
	  PORT MAP ( 
		arctan => wire_cata_0_cordic_atan_arctan,
		indexbit => indexbitff(0)
	  );
	cata_10_cordic_atan :  coshw_altfp_sincos_cordic_atan_k6b
	  PORT MAP ( 
		arctan => wire_cata_10_cordic_atan_arctan,
		indexbit => indexbitff(10)
	  );
	cata_11_cordic_atan :  coshw_altfp_sincos_cordic_atan_l6b
	  PORT MAP ( 
		arctan => wire_cata_11_cordic_atan_arctan,
		indexbit => indexbitff(11)
	  );
	cata_12_cordic_atan :  coshw_altfp_sincos_cordic_atan_m6b
	  PORT MAP ( 
		arctan => wire_cata_12_cordic_atan_arctan,
		indexbit => indexbitff(12)
	  );
	cata_13_cordic_atan :  coshw_altfp_sincos_cordic_atan_n6b
	  PORT MAP ( 
		arctan => wire_cata_13_cordic_atan_arctan,
		indexbit => indexbitff(13)
	  );
	cata_1_cordic_atan :  coshw_altfp_sincos_cordic_atan_45b
	  PORT MAP ( 
		arctan => wire_cata_1_cordic_atan_arctan,
		indexbit => indexbitff(1)
	  );
	cata_2_cordic_atan :  coshw_altfp_sincos_cordic_atan_55b
	  PORT MAP ( 
		arctan => wire_cata_2_cordic_atan_arctan,
		indexbit => indexbitff(2)
	  );
	cata_3_cordic_atan :  coshw_altfp_sincos_cordic_atan_65b
	  PORT MAP ( 
		arctan => wire_cata_3_cordic_atan_arctan,
		indexbit => indexbitff(3)
	  );
	cata_4_cordic_atan :  coshw_altfp_sincos_cordic_atan_75b
	  PORT MAP ( 
		arctan => wire_cata_4_cordic_atan_arctan,
		indexbit => indexbitff(4)
	  );
	cata_5_cordic_atan :  coshw_altfp_sincos_cordic_atan_85b
	  PORT MAP ( 
		arctan => wire_cata_5_cordic_atan_arctan,
		indexbit => indexbitff(5)
	  );
	cata_6_cordic_atan :  coshw_altfp_sincos_cordic_atan_95b
	  PORT MAP ( 
		arctan => wire_cata_6_cordic_atan_arctan,
		indexbit => indexbitff(6)
	  );
	cata_7_cordic_atan :  coshw_altfp_sincos_cordic_atan_a5b
	  PORT MAP ( 
		arctan => wire_cata_7_cordic_atan_arctan,
		indexbit => indexbitff(7)
	  );
	cata_8_cordic_atan :  coshw_altfp_sincos_cordic_atan_b5b
	  PORT MAP ( 
		arctan => wire_cata_8_cordic_atan_arctan,
		indexbit => indexbitff(8)
	  );
	cata_9_cordic_atan :  coshw_altfp_sincos_cordic_atan_c5b
	  PORT MAP ( 
		arctan => wire_cata_9_cordic_atan_arctan,
		indexbit => indexbitff(9)
	  );
	cxs :  coshw_altfp_sincos_cordic_start_509
	  PORT MAP ( 
		index => startindex_w,
		value => wire_cxs_value
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cdaff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cdaff_0 <= delay_input_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cdaff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cdaff_1 <= cdaff_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cdaff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cdaff_2 <= cdaff_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN indexbitff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN indexbitff <= ( indexbitff(15 DOWNTO 0) & indexbit);
			END IF;
		END IF;
	END PROCESS;
	wire_indexbitff_w_lg_w_q_range448w546w(0) <= NOT wire_indexbitff_w_q_range448w(0);
	wire_indexbitff_w_lg_w_q_range477w7967w(0) <= NOT wire_indexbitff_w_q_range477w(0);
	wire_indexbitff_w_lg_w_q_range480w8718w(0) <= NOT wire_indexbitff_w_q_range480w(0);
	wire_indexbitff_w_lg_w_q_range483w9464w(0) <= NOT wire_indexbitff_w_q_range483w(0);
	wire_indexbitff_w_lg_w_q_range9992w9995w(0) <= NOT wire_indexbitff_w_q_range9992w(0);
	wire_indexbitff_w_lg_w_q_range450w983w(0) <= NOT wire_indexbitff_w_q_range450w(0);
	wire_indexbitff_w_lg_w_q_range453w1779w(0) <= NOT wire_indexbitff_w_q_range453w(0);
	wire_indexbitff_w_lg_w_q_range456w2570w(0) <= NOT wire_indexbitff_w_q_range456w(0);
	wire_indexbitff_w_lg_w_q_range459w3356w(0) <= NOT wire_indexbitff_w_q_range459w(0);
	wire_indexbitff_w_lg_w_q_range462w4137w(0) <= NOT wire_indexbitff_w_q_range462w(0);
	wire_indexbitff_w_lg_w_q_range465w4913w(0) <= NOT wire_indexbitff_w_q_range465w(0);
	wire_indexbitff_w_lg_w_q_range468w5684w(0) <= NOT wire_indexbitff_w_q_range468w(0);
	wire_indexbitff_w_lg_w_q_range471w6450w(0) <= NOT wire_indexbitff_w_q_range471w(0);
	wire_indexbitff_w_lg_w_q_range474w7211w(0) <= NOT wire_indexbitff_w_q_range474w(0);
	wire_indexbitff_w_q_range448w(0) <= indexbitff(0);
	wire_indexbitff_w_q_range477w(0) <= indexbitff(10);
	wire_indexbitff_w_q_range480w(0) <= indexbitff(11);
	wire_indexbitff_w_q_range483w(0) <= indexbitff(12);
	wire_indexbitff_w_q_range9992w(0) <= indexbitff(16);
	wire_indexbitff_w_q_range450w(0) <= indexbitff(1);
	wire_indexbitff_w_q_range453w(0) <= indexbitff(2);
	wire_indexbitff_w_q_range456w(0) <= indexbitff(3);
	wire_indexbitff_w_q_range459w(0) <= indexbitff(4);
	wire_indexbitff_w_q_range462w(0) <= indexbitff(5);
	wire_indexbitff_w_q_range465w(0) <= indexbitff(6);
	wire_indexbitff_w_q_range468w(0) <= indexbitff(7);
	wire_indexbitff_w_q_range471w(0) <= indexbitff(8);
	wire_indexbitff_w_q_range474w(0) <= indexbitff(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sincosbitff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN sincosbitff <= ( sincosbitff(15 DOWNTO 0) & sincosbit);
			END IF;
		END IF;
	END PROCESS;
	wire_sincosbitff_w_lg_w_q_range535w9982w(0) <= NOT wire_sincosbitff_w_q_range535w(0);
	wire_sincosbitff_w_lg_w_q_range9989w9990w(0) <= NOT wire_sincosbitff_w_q_range9989w(0);
	wire_sincosbitff_w_q_range535w(0) <= sincosbitff(13);
	wire_sincosbitff_w_q_range9989w(0) <= sincosbitff(16);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sincosff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN sincosff <= wire_sincos_add_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_0 <= x_start_node_w;
			END IF;
		END IF;
	END PROCESS;
	wire_x_pipeff_0_w_lg_w_q_range547w548w(0) <= wire_x_pipeff_0_w_q_range547w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range584w601w(0) <= wire_x_pipeff_0_w_q_range584w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range584w585w(0) <= wire_x_pipeff_0_w_q_range584w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range589w606w(0) <= wire_x_pipeff_0_w_q_range589w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range589w590w(0) <= wire_x_pipeff_0_w_q_range589w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range594w611w(0) <= wire_x_pipeff_0_w_q_range594w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range594w595w(0) <= wire_x_pipeff_0_w_q_range594w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range599w616w(0) <= wire_x_pipeff_0_w_q_range599w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range599w600w(0) <= wire_x_pipeff_0_w_q_range599w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range604w621w(0) <= wire_x_pipeff_0_w_q_range604w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range604w605w(0) <= wire_x_pipeff_0_w_q_range604w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range609w626w(0) <= wire_x_pipeff_0_w_q_range609w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range609w610w(0) <= wire_x_pipeff_0_w_q_range609w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range614w631w(0) <= wire_x_pipeff_0_w_q_range614w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range614w615w(0) <= wire_x_pipeff_0_w_q_range614w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range619w636w(0) <= wire_x_pipeff_0_w_q_range619w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range619w620w(0) <= wire_x_pipeff_0_w_q_range619w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range624w641w(0) <= wire_x_pipeff_0_w_q_range624w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range624w625w(0) <= wire_x_pipeff_0_w_q_range624w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range629w646w(0) <= wire_x_pipeff_0_w_q_range629w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range629w630w(0) <= wire_x_pipeff_0_w_q_range629w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range554w555w(0) <= wire_x_pipeff_0_w_q_range554w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range634w651w(0) <= wire_x_pipeff_0_w_q_range634w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range634w635w(0) <= wire_x_pipeff_0_w_q_range634w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range639w656w(0) <= wire_x_pipeff_0_w_q_range639w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range639w640w(0) <= wire_x_pipeff_0_w_q_range639w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range644w661w(0) <= wire_x_pipeff_0_w_q_range644w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range644w645w(0) <= wire_x_pipeff_0_w_q_range644w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range649w666w(0) <= wire_x_pipeff_0_w_q_range649w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range649w650w(0) <= wire_x_pipeff_0_w_q_range649w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range654w671w(0) <= wire_x_pipeff_0_w_q_range654w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range654w655w(0) <= wire_x_pipeff_0_w_q_range654w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range659w676w(0) <= wire_x_pipeff_0_w_q_range659w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range659w660w(0) <= wire_x_pipeff_0_w_q_range659w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range664w681w(0) <= wire_x_pipeff_0_w_q_range664w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range664w665w(0) <= wire_x_pipeff_0_w_q_range664w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range669w686w(0) <= wire_x_pipeff_0_w_q_range669w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range669w670w(0) <= wire_x_pipeff_0_w_q_range669w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range674w691w(0) <= wire_x_pipeff_0_w_q_range674w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range674w675w(0) <= wire_x_pipeff_0_w_q_range674w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range679w694w(0) <= wire_x_pipeff_0_w_q_range679w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range679w680w(0) <= wire_x_pipeff_0_w_q_range679w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range560w561w(0) <= wire_x_pipeff_0_w_q_range560w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range684w696w(0) <= wire_x_pipeff_0_w_q_range684w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range684w685w(0) <= wire_x_pipeff_0_w_q_range684w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range689w690w(0) <= wire_x_pipeff_0_w_q_range689w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range544w566w(0) <= wire_x_pipeff_0_w_q_range544w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range544w545w(0) <= wire_x_pipeff_0_w_q_range544w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range552w571w(0) <= wire_x_pipeff_0_w_q_range552w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range552w553w(0) <= wire_x_pipeff_0_w_q_range552w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range558w576w(0) <= wire_x_pipeff_0_w_q_range558w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range558w559w(0) <= wire_x_pipeff_0_w_q_range558w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range564w581w(0) <= wire_x_pipeff_0_w_q_range564w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range564w565w(0) <= wire_x_pipeff_0_w_q_range564w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range569w586w(0) <= wire_x_pipeff_0_w_q_range569w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range569w570w(0) <= wire_x_pipeff_0_w_q_range569w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range574w591w(0) <= wire_x_pipeff_0_w_q_range574w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range574w575w(0) <= wire_x_pipeff_0_w_q_range574w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range579w596w(0) <= wire_x_pipeff_0_w_q_range579w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_q_range579w580w(0) <= wire_x_pipeff_0_w_q_range579w(0) AND wire_indexbitff_w_q_range448w(0);
	wire_x_pipeff_0_w_lg_w_q_range689w698w(0) <= wire_x_pipeff_0_w_q_range689w(0) AND wire_indexbitff_w_lg_w_q_range448w546w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range547w548w549w(0) <= wire_x_pipeff_0_w_lg_w_q_range547w548w(0) OR wire_x_pipeff_0_w_lg_w_q_range544w545w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range584w601w602w(0) <= wire_x_pipeff_0_w_lg_w_q_range584w601w(0) OR wire_x_pipeff_0_w_lg_w_q_range599w600w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range589w606w607w(0) <= wire_x_pipeff_0_w_lg_w_q_range589w606w(0) OR wire_x_pipeff_0_w_lg_w_q_range604w605w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range594w611w612w(0) <= wire_x_pipeff_0_w_lg_w_q_range594w611w(0) OR wire_x_pipeff_0_w_lg_w_q_range609w610w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range599w616w617w(0) <= wire_x_pipeff_0_w_lg_w_q_range599w616w(0) OR wire_x_pipeff_0_w_lg_w_q_range614w615w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range604w621w622w(0) <= wire_x_pipeff_0_w_lg_w_q_range604w621w(0) OR wire_x_pipeff_0_w_lg_w_q_range619w620w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range609w626w627w(0) <= wire_x_pipeff_0_w_lg_w_q_range609w626w(0) OR wire_x_pipeff_0_w_lg_w_q_range624w625w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range614w631w632w(0) <= wire_x_pipeff_0_w_lg_w_q_range614w631w(0) OR wire_x_pipeff_0_w_lg_w_q_range629w630w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range619w636w637w(0) <= wire_x_pipeff_0_w_lg_w_q_range619w636w(0) OR wire_x_pipeff_0_w_lg_w_q_range634w635w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range624w641w642w(0) <= wire_x_pipeff_0_w_lg_w_q_range624w641w(0) OR wire_x_pipeff_0_w_lg_w_q_range639w640w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range629w646w647w(0) <= wire_x_pipeff_0_w_lg_w_q_range629w646w(0) OR wire_x_pipeff_0_w_lg_w_q_range644w645w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range554w555w556w(0) <= wire_x_pipeff_0_w_lg_w_q_range554w555w(0) OR wire_x_pipeff_0_w_lg_w_q_range552w553w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range634w651w652w(0) <= wire_x_pipeff_0_w_lg_w_q_range634w651w(0) OR wire_x_pipeff_0_w_lg_w_q_range649w650w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range639w656w657w(0) <= wire_x_pipeff_0_w_lg_w_q_range639w656w(0) OR wire_x_pipeff_0_w_lg_w_q_range654w655w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range644w661w662w(0) <= wire_x_pipeff_0_w_lg_w_q_range644w661w(0) OR wire_x_pipeff_0_w_lg_w_q_range659w660w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range649w666w667w(0) <= wire_x_pipeff_0_w_lg_w_q_range649w666w(0) OR wire_x_pipeff_0_w_lg_w_q_range664w665w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range654w671w672w(0) <= wire_x_pipeff_0_w_lg_w_q_range654w671w(0) OR wire_x_pipeff_0_w_lg_w_q_range669w670w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range659w676w677w(0) <= wire_x_pipeff_0_w_lg_w_q_range659w676w(0) OR wire_x_pipeff_0_w_lg_w_q_range674w675w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range664w681w682w(0) <= wire_x_pipeff_0_w_lg_w_q_range664w681w(0) OR wire_x_pipeff_0_w_lg_w_q_range679w680w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range669w686w687w(0) <= wire_x_pipeff_0_w_lg_w_q_range669w686w(0) OR wire_x_pipeff_0_w_lg_w_q_range684w685w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range674w691w692w(0) <= wire_x_pipeff_0_w_lg_w_q_range674w691w(0) OR wire_x_pipeff_0_w_lg_w_q_range689w690w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range560w561w562w(0) <= wire_x_pipeff_0_w_lg_w_q_range560w561w(0) OR wire_x_pipeff_0_w_lg_w_q_range558w559w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range544w566w567w(0) <= wire_x_pipeff_0_w_lg_w_q_range544w566w(0) OR wire_x_pipeff_0_w_lg_w_q_range564w565w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range552w571w572w(0) <= wire_x_pipeff_0_w_lg_w_q_range552w571w(0) OR wire_x_pipeff_0_w_lg_w_q_range569w570w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range558w576w577w(0) <= wire_x_pipeff_0_w_lg_w_q_range558w576w(0) OR wire_x_pipeff_0_w_lg_w_q_range574w575w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range564w581w582w(0) <= wire_x_pipeff_0_w_lg_w_q_range564w581w(0) OR wire_x_pipeff_0_w_lg_w_q_range579w580w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range569w586w587w(0) <= wire_x_pipeff_0_w_lg_w_q_range569w586w(0) OR wire_x_pipeff_0_w_lg_w_q_range584w585w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range574w591w592w(0) <= wire_x_pipeff_0_w_lg_w_q_range574w591w(0) OR wire_x_pipeff_0_w_lg_w_q_range589w590w(0);
	wire_x_pipeff_0_w_lg_w_lg_w_q_range579w596w597w(0) <= wire_x_pipeff_0_w_lg_w_q_range579w596w(0) OR wire_x_pipeff_0_w_lg_w_q_range594w595w(0);
	wire_x_pipeff_0_w_q_range547w(0) <= x_pipeff_0(0);
	wire_x_pipeff_0_w_q_range584w(0) <= x_pipeff_0(10);
	wire_x_pipeff_0_w_q_range589w(0) <= x_pipeff_0(11);
	wire_x_pipeff_0_w_q_range594w(0) <= x_pipeff_0(12);
	wire_x_pipeff_0_w_q_range599w(0) <= x_pipeff_0(13);
	wire_x_pipeff_0_w_q_range604w(0) <= x_pipeff_0(14);
	wire_x_pipeff_0_w_q_range609w(0) <= x_pipeff_0(15);
	wire_x_pipeff_0_w_q_range614w(0) <= x_pipeff_0(16);
	wire_x_pipeff_0_w_q_range619w(0) <= x_pipeff_0(17);
	wire_x_pipeff_0_w_q_range624w(0) <= x_pipeff_0(18);
	wire_x_pipeff_0_w_q_range629w(0) <= x_pipeff_0(19);
	wire_x_pipeff_0_w_q_range554w(0) <= x_pipeff_0(1);
	wire_x_pipeff_0_w_q_range634w(0) <= x_pipeff_0(20);
	wire_x_pipeff_0_w_q_range639w(0) <= x_pipeff_0(21);
	wire_x_pipeff_0_w_q_range644w(0) <= x_pipeff_0(22);
	wire_x_pipeff_0_w_q_range649w(0) <= x_pipeff_0(23);
	wire_x_pipeff_0_w_q_range654w(0) <= x_pipeff_0(24);
	wire_x_pipeff_0_w_q_range659w(0) <= x_pipeff_0(25);
	wire_x_pipeff_0_w_q_range664w(0) <= x_pipeff_0(26);
	wire_x_pipeff_0_w_q_range669w(0) <= x_pipeff_0(27);
	wire_x_pipeff_0_w_q_range674w(0) <= x_pipeff_0(28);
	wire_x_pipeff_0_w_q_range679w(0) <= x_pipeff_0(29);
	wire_x_pipeff_0_w_q_range560w(0) <= x_pipeff_0(2);
	wire_x_pipeff_0_w_q_range684w(0) <= x_pipeff_0(30);
	wire_x_pipeff_0_w_q_range689w(0) <= x_pipeff_0(31);
	wire_x_pipeff_0_w_q_range544w(0) <= x_pipeff_0(3);
	wire_x_pipeff_0_w_q_range552w(0) <= x_pipeff_0(4);
	wire_x_pipeff_0_w_q_range558w(0) <= x_pipeff_0(5);
	wire_x_pipeff_0_w_q_range564w(0) <= x_pipeff_0(6);
	wire_x_pipeff_0_w_q_range569w(0) <= x_pipeff_0(7);
	wire_x_pipeff_0_w_q_range574w(0) <= x_pipeff_0(8);
	wire_x_pipeff_0_w_q_range579w(0) <= x_pipeff_0(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_1 <= x_pipeff_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_10 <= x_pipenode_10_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_11 <= x_pipenode_11_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_12 <= x_pipenode_12_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_13 <= x_pipenode_13_w;
			END IF;
		END IF;
	END PROCESS;
	loop32 : FOR i IN 0 TO 31 GENERATE 
		wire_x_pipeff_13_w_lg_q9987w(i) <= x_pipeff_13(i) AND wire_sincosbitff_w_lg_w_q_range535w9982w(0);
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 31 GENERATE 
		wire_x_pipeff_13_w_lg_q9984w(i) <= x_pipeff_13(i) AND wire_sincosbitff_w_q_range535w(0);
	END GENERATE loop33;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_2 <= x_pipenode_2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_3 <= x_pipenode_3_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_4 <= x_pipenode_4_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_5 <= x_pipenode_5_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_6 <= x_pipenode_6_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_7 <= x_pipenode_7_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_8 <= x_pipenode_8_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN x_pipeff_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN x_pipeff_9 <= x_pipenode_9_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(0) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(0) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(1) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(1) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(2) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(2) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(3) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(3) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(4) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(4) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(5) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(5) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(6) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(6) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(7) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(7) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(8) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(8) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(9) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(9) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(10) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(10) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(11) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(11) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(12) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(12) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(13) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(13) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(14) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(14) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(15) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(15) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(16) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(16) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(17) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(17) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(18) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(18) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(19) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(19) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(20) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(20) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(21) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(21) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(22) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(22) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(23) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(23) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(24) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(24) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(25) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(25) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(26) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(26) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(27) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(27) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(28) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(28) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(29) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(29) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(30) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(30) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_0(31) <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_0(31) <= '0';
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_1 <= wire_y_pipeff1_add_result;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_1_w_lg_w_q_range770w771w(0) <= NOT wire_y_pipeff_1_w_q_range770w(0);
	wire_y_pipeff_1_w_lg_w_q_range776w777w(0) <= NOT wire_y_pipeff_1_w_q_range776w(0);
	wire_y_pipeff_1_w_lg_w_q_range782w783w(0) <= NOT wire_y_pipeff_1_w_q_range782w(0);
	wire_y_pipeff_1_w_lg_w_q_range788w789w(0) <= NOT wire_y_pipeff_1_w_q_range788w(0);
	wire_y_pipeff_1_w_lg_w_q_range794w795w(0) <= NOT wire_y_pipeff_1_w_q_range794w(0);
	wire_y_pipeff_1_w_lg_w_q_range800w801w(0) <= NOT wire_y_pipeff_1_w_q_range800w(0);
	wire_y_pipeff_1_w_lg_w_q_range806w807w(0) <= NOT wire_y_pipeff_1_w_q_range806w(0);
	wire_y_pipeff_1_w_lg_w_q_range812w813w(0) <= NOT wire_y_pipeff_1_w_q_range812w(0);
	wire_y_pipeff_1_w_lg_w_q_range818w819w(0) <= NOT wire_y_pipeff_1_w_q_range818w(0);
	wire_y_pipeff_1_w_lg_w_q_range824w825w(0) <= NOT wire_y_pipeff_1_w_q_range824w(0);
	wire_y_pipeff_1_w_lg_w_q_range717w718w(0) <= NOT wire_y_pipeff_1_w_q_range717w(0);
	wire_y_pipeff_1_w_lg_w_q_range830w831w(0) <= NOT wire_y_pipeff_1_w_q_range830w(0);
	wire_y_pipeff_1_w_lg_w_q_range836w837w(0) <= NOT wire_y_pipeff_1_w_q_range836w(0);
	wire_y_pipeff_1_w_lg_w_q_range842w843w(0) <= NOT wire_y_pipeff_1_w_q_range842w(0);
	wire_y_pipeff_1_w_lg_w_q_range848w849w(0) <= NOT wire_y_pipeff_1_w_q_range848w(0);
	wire_y_pipeff_1_w_lg_w_q_range854w855w(0) <= NOT wire_y_pipeff_1_w_q_range854w(0);
	wire_y_pipeff_1_w_lg_w_q_range860w861w(0) <= NOT wire_y_pipeff_1_w_q_range860w(0);
	wire_y_pipeff_1_w_lg_w_q_range866w867w(0) <= NOT wire_y_pipeff_1_w_q_range866w(0);
	wire_y_pipeff_1_w_lg_w_q_range872w873w(0) <= NOT wire_y_pipeff_1_w_q_range872w(0);
	wire_y_pipeff_1_w_lg_w_q_range878w879w(0) <= NOT wire_y_pipeff_1_w_q_range878w(0);
	wire_y_pipeff_1_w_lg_w_q_range884w885w(0) <= NOT wire_y_pipeff_1_w_q_range884w(0);
	wire_y_pipeff_1_w_lg_w_q_range722w723w(0) <= NOT wire_y_pipeff_1_w_q_range722w(0);
	wire_y_pipeff_1_w_lg_w_q_range890w891w(0) <= NOT wire_y_pipeff_1_w_q_range890w(0);
	wire_y_pipeff_1_w_lg_w_q_range700w701w(0) <= NOT wire_y_pipeff_1_w_q_range700w(0);
	wire_y_pipeff_1_w_lg_w_q_range728w729w(0) <= NOT wire_y_pipeff_1_w_q_range728w(0);
	wire_y_pipeff_1_w_lg_w_q_range734w735w(0) <= NOT wire_y_pipeff_1_w_q_range734w(0);
	wire_y_pipeff_1_w_lg_w_q_range740w741w(0) <= NOT wire_y_pipeff_1_w_q_range740w(0);
	wire_y_pipeff_1_w_lg_w_q_range746w747w(0) <= NOT wire_y_pipeff_1_w_q_range746w(0);
	wire_y_pipeff_1_w_lg_w_q_range752w753w(0) <= NOT wire_y_pipeff_1_w_q_range752w(0);
	wire_y_pipeff_1_w_lg_w_q_range758w759w(0) <= NOT wire_y_pipeff_1_w_q_range758w(0);
	wire_y_pipeff_1_w_lg_w_q_range764w765w(0) <= NOT wire_y_pipeff_1_w_q_range764w(0);
	wire_y_pipeff_1_w_q_range770w(0) <= y_pipeff_1(10);
	wire_y_pipeff_1_w_q_range776w(0) <= y_pipeff_1(11);
	wire_y_pipeff_1_w_q_range782w(0) <= y_pipeff_1(12);
	wire_y_pipeff_1_w_q_range788w(0) <= y_pipeff_1(13);
	wire_y_pipeff_1_w_q_range794w(0) <= y_pipeff_1(14);
	wire_y_pipeff_1_w_q_range800w(0) <= y_pipeff_1(15);
	wire_y_pipeff_1_w_q_range806w(0) <= y_pipeff_1(16);
	wire_y_pipeff_1_w_q_range812w(0) <= y_pipeff_1(17);
	wire_y_pipeff_1_w_q_range818w(0) <= y_pipeff_1(18);
	wire_y_pipeff_1_w_q_range824w(0) <= y_pipeff_1(19);
	wire_y_pipeff_1_w_q_range717w(0) <= y_pipeff_1(1);
	wire_y_pipeff_1_w_q_range830w(0) <= y_pipeff_1(20);
	wire_y_pipeff_1_w_q_range836w(0) <= y_pipeff_1(21);
	wire_y_pipeff_1_w_q_range842w(0) <= y_pipeff_1(22);
	wire_y_pipeff_1_w_q_range848w(0) <= y_pipeff_1(23);
	wire_y_pipeff_1_w_q_range854w(0) <= y_pipeff_1(24);
	wire_y_pipeff_1_w_q_range860w(0) <= y_pipeff_1(25);
	wire_y_pipeff_1_w_q_range866w(0) <= y_pipeff_1(26);
	wire_y_pipeff_1_w_q_range872w(0) <= y_pipeff_1(27);
	wire_y_pipeff_1_w_q_range878w(0) <= y_pipeff_1(28);
	wire_y_pipeff_1_w_q_range884w(0) <= y_pipeff_1(29);
	wire_y_pipeff_1_w_q_range722w(0) <= y_pipeff_1(2);
	wire_y_pipeff_1_w_q_range890w(0) <= y_pipeff_1(30);
	wire_y_pipeff_1_w_q_range700w(0) <= y_pipeff_1(31);
	wire_y_pipeff_1_w_q_range728w(0) <= y_pipeff_1(3);
	wire_y_pipeff_1_w_q_range734w(0) <= y_pipeff_1(4);
	wire_y_pipeff_1_w_q_range740w(0) <= y_pipeff_1(5);
	wire_y_pipeff_1_w_q_range746w(0) <= y_pipeff_1(6);
	wire_y_pipeff_1_w_q_range752w(0) <= y_pipeff_1(7);
	wire_y_pipeff_1_w_q_range758w(0) <= y_pipeff_1(8);
	wire_y_pipeff_1_w_q_range764w(0) <= y_pipeff_1(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_10 <= y_pipenode_10_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_10_w_lg_w_q_range7782w7783w(0) <= NOT wire_y_pipeff_10_w_q_range7782w(0);
	wire_y_pipeff_10_w_lg_w_q_range7787w7788w(0) <= NOT wire_y_pipeff_10_w_q_range7787w(0);
	wire_y_pipeff_10_w_lg_w_q_range7793w7794w(0) <= NOT wire_y_pipeff_10_w_q_range7793w(0);
	wire_y_pipeff_10_w_lg_w_q_range7799w7800w(0) <= NOT wire_y_pipeff_10_w_q_range7799w(0);
	wire_y_pipeff_10_w_lg_w_q_range7805w7806w(0) <= NOT wire_y_pipeff_10_w_q_range7805w(0);
	wire_y_pipeff_10_w_lg_w_q_range7811w7812w(0) <= NOT wire_y_pipeff_10_w_q_range7811w(0);
	wire_y_pipeff_10_w_lg_w_q_range7817w7818w(0) <= NOT wire_y_pipeff_10_w_q_range7817w(0);
	wire_y_pipeff_10_w_lg_w_q_range7823w7824w(0) <= NOT wire_y_pipeff_10_w_q_range7823w(0);
	wire_y_pipeff_10_w_lg_w_q_range7829w7830w(0) <= NOT wire_y_pipeff_10_w_q_range7829w(0);
	wire_y_pipeff_10_w_lg_w_q_range7835w7836w(0) <= NOT wire_y_pipeff_10_w_q_range7835w(0);
	wire_y_pipeff_10_w_lg_w_q_range7841w7842w(0) <= NOT wire_y_pipeff_10_w_q_range7841w(0);
	wire_y_pipeff_10_w_lg_w_q_range7847w7848w(0) <= NOT wire_y_pipeff_10_w_q_range7847w(0);
	wire_y_pipeff_10_w_lg_w_q_range7853w7854w(0) <= NOT wire_y_pipeff_10_w_q_range7853w(0);
	wire_y_pipeff_10_w_lg_w_q_range7859w7860w(0) <= NOT wire_y_pipeff_10_w_q_range7859w(0);
	wire_y_pipeff_10_w_lg_w_q_range7865w7866w(0) <= NOT wire_y_pipeff_10_w_q_range7865w(0);
	wire_y_pipeff_10_w_lg_w_q_range7871w7872w(0) <= NOT wire_y_pipeff_10_w_q_range7871w(0);
	wire_y_pipeff_10_w_lg_w_q_range7877w7878w(0) <= NOT wire_y_pipeff_10_w_q_range7877w(0);
	wire_y_pipeff_10_w_lg_w_q_range7883w7884w(0) <= NOT wire_y_pipeff_10_w_q_range7883w(0);
	wire_y_pipeff_10_w_lg_w_q_range7889w7890w(0) <= NOT wire_y_pipeff_10_w_q_range7889w(0);
	wire_y_pipeff_10_w_lg_w_q_range7895w7896w(0) <= NOT wire_y_pipeff_10_w_q_range7895w(0);
	wire_y_pipeff_10_w_lg_w_q_range7901w7902w(0) <= NOT wire_y_pipeff_10_w_q_range7901w(0);
	wire_y_pipeff_10_w_lg_w_q_range7729w7730w(0) <= NOT wire_y_pipeff_10_w_q_range7729w(0);
	wire_y_pipeff_10_w_q_range7782w(0) <= y_pipeff_10(10);
	wire_y_pipeff_10_w_q_range7787w(0) <= y_pipeff_10(11);
	wire_y_pipeff_10_w_q_range7793w(0) <= y_pipeff_10(12);
	wire_y_pipeff_10_w_q_range7799w(0) <= y_pipeff_10(13);
	wire_y_pipeff_10_w_q_range7805w(0) <= y_pipeff_10(14);
	wire_y_pipeff_10_w_q_range7811w(0) <= y_pipeff_10(15);
	wire_y_pipeff_10_w_q_range7817w(0) <= y_pipeff_10(16);
	wire_y_pipeff_10_w_q_range7823w(0) <= y_pipeff_10(17);
	wire_y_pipeff_10_w_q_range7829w(0) <= y_pipeff_10(18);
	wire_y_pipeff_10_w_q_range7835w(0) <= y_pipeff_10(19);
	wire_y_pipeff_10_w_q_range7841w(0) <= y_pipeff_10(20);
	wire_y_pipeff_10_w_q_range7847w(0) <= y_pipeff_10(21);
	wire_y_pipeff_10_w_q_range7853w(0) <= y_pipeff_10(22);
	wire_y_pipeff_10_w_q_range7859w(0) <= y_pipeff_10(23);
	wire_y_pipeff_10_w_q_range7865w(0) <= y_pipeff_10(24);
	wire_y_pipeff_10_w_q_range7871w(0) <= y_pipeff_10(25);
	wire_y_pipeff_10_w_q_range7877w(0) <= y_pipeff_10(26);
	wire_y_pipeff_10_w_q_range7883w(0) <= y_pipeff_10(27);
	wire_y_pipeff_10_w_q_range7889w(0) <= y_pipeff_10(28);
	wire_y_pipeff_10_w_q_range7895w(0) <= y_pipeff_10(29);
	wire_y_pipeff_10_w_q_range7901w(0) <= y_pipeff_10(30);
	wire_y_pipeff_10_w_q_range7729w(0) <= y_pipeff_10(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_11 <= y_pipenode_11_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_11_w_lg_w_q_range8542w8543w(0) <= NOT wire_y_pipeff_11_w_q_range8542w(0);
	wire_y_pipeff_11_w_lg_w_q_range8547w8548w(0) <= NOT wire_y_pipeff_11_w_q_range8547w(0);
	wire_y_pipeff_11_w_lg_w_q_range8553w8554w(0) <= NOT wire_y_pipeff_11_w_q_range8553w(0);
	wire_y_pipeff_11_w_lg_w_q_range8559w8560w(0) <= NOT wire_y_pipeff_11_w_q_range8559w(0);
	wire_y_pipeff_11_w_lg_w_q_range8565w8566w(0) <= NOT wire_y_pipeff_11_w_q_range8565w(0);
	wire_y_pipeff_11_w_lg_w_q_range8571w8572w(0) <= NOT wire_y_pipeff_11_w_q_range8571w(0);
	wire_y_pipeff_11_w_lg_w_q_range8577w8578w(0) <= NOT wire_y_pipeff_11_w_q_range8577w(0);
	wire_y_pipeff_11_w_lg_w_q_range8583w8584w(0) <= NOT wire_y_pipeff_11_w_q_range8583w(0);
	wire_y_pipeff_11_w_lg_w_q_range8589w8590w(0) <= NOT wire_y_pipeff_11_w_q_range8589w(0);
	wire_y_pipeff_11_w_lg_w_q_range8595w8596w(0) <= NOT wire_y_pipeff_11_w_q_range8595w(0);
	wire_y_pipeff_11_w_lg_w_q_range8601w8602w(0) <= NOT wire_y_pipeff_11_w_q_range8601w(0);
	wire_y_pipeff_11_w_lg_w_q_range8607w8608w(0) <= NOT wire_y_pipeff_11_w_q_range8607w(0);
	wire_y_pipeff_11_w_lg_w_q_range8613w8614w(0) <= NOT wire_y_pipeff_11_w_q_range8613w(0);
	wire_y_pipeff_11_w_lg_w_q_range8619w8620w(0) <= NOT wire_y_pipeff_11_w_q_range8619w(0);
	wire_y_pipeff_11_w_lg_w_q_range8625w8626w(0) <= NOT wire_y_pipeff_11_w_q_range8625w(0);
	wire_y_pipeff_11_w_lg_w_q_range8631w8632w(0) <= NOT wire_y_pipeff_11_w_q_range8631w(0);
	wire_y_pipeff_11_w_lg_w_q_range8637w8638w(0) <= NOT wire_y_pipeff_11_w_q_range8637w(0);
	wire_y_pipeff_11_w_lg_w_q_range8643w8644w(0) <= NOT wire_y_pipeff_11_w_q_range8643w(0);
	wire_y_pipeff_11_w_lg_w_q_range8649w8650w(0) <= NOT wire_y_pipeff_11_w_q_range8649w(0);
	wire_y_pipeff_11_w_lg_w_q_range8655w8656w(0) <= NOT wire_y_pipeff_11_w_q_range8655w(0);
	wire_y_pipeff_11_w_lg_w_q_range8485w8486w(0) <= NOT wire_y_pipeff_11_w_q_range8485w(0);
	wire_y_pipeff_11_w_q_range8542w(0) <= y_pipeff_11(11);
	wire_y_pipeff_11_w_q_range8547w(0) <= y_pipeff_11(12);
	wire_y_pipeff_11_w_q_range8553w(0) <= y_pipeff_11(13);
	wire_y_pipeff_11_w_q_range8559w(0) <= y_pipeff_11(14);
	wire_y_pipeff_11_w_q_range8565w(0) <= y_pipeff_11(15);
	wire_y_pipeff_11_w_q_range8571w(0) <= y_pipeff_11(16);
	wire_y_pipeff_11_w_q_range8577w(0) <= y_pipeff_11(17);
	wire_y_pipeff_11_w_q_range8583w(0) <= y_pipeff_11(18);
	wire_y_pipeff_11_w_q_range8589w(0) <= y_pipeff_11(19);
	wire_y_pipeff_11_w_q_range8595w(0) <= y_pipeff_11(20);
	wire_y_pipeff_11_w_q_range8601w(0) <= y_pipeff_11(21);
	wire_y_pipeff_11_w_q_range8607w(0) <= y_pipeff_11(22);
	wire_y_pipeff_11_w_q_range8613w(0) <= y_pipeff_11(23);
	wire_y_pipeff_11_w_q_range8619w(0) <= y_pipeff_11(24);
	wire_y_pipeff_11_w_q_range8625w(0) <= y_pipeff_11(25);
	wire_y_pipeff_11_w_q_range8631w(0) <= y_pipeff_11(26);
	wire_y_pipeff_11_w_q_range8637w(0) <= y_pipeff_11(27);
	wire_y_pipeff_11_w_q_range8643w(0) <= y_pipeff_11(28);
	wire_y_pipeff_11_w_q_range8649w(0) <= y_pipeff_11(29);
	wire_y_pipeff_11_w_q_range8655w(0) <= y_pipeff_11(30);
	wire_y_pipeff_11_w_q_range8485w(0) <= y_pipeff_11(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_12 <= y_pipenode_12_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_12_w_lg_w_q_range9297w9298w(0) <= NOT wire_y_pipeff_12_w_q_range9297w(0);
	wire_y_pipeff_12_w_lg_w_q_range9302w9303w(0) <= NOT wire_y_pipeff_12_w_q_range9302w(0);
	wire_y_pipeff_12_w_lg_w_q_range9308w9309w(0) <= NOT wire_y_pipeff_12_w_q_range9308w(0);
	wire_y_pipeff_12_w_lg_w_q_range9314w9315w(0) <= NOT wire_y_pipeff_12_w_q_range9314w(0);
	wire_y_pipeff_12_w_lg_w_q_range9320w9321w(0) <= NOT wire_y_pipeff_12_w_q_range9320w(0);
	wire_y_pipeff_12_w_lg_w_q_range9326w9327w(0) <= NOT wire_y_pipeff_12_w_q_range9326w(0);
	wire_y_pipeff_12_w_lg_w_q_range9332w9333w(0) <= NOT wire_y_pipeff_12_w_q_range9332w(0);
	wire_y_pipeff_12_w_lg_w_q_range9338w9339w(0) <= NOT wire_y_pipeff_12_w_q_range9338w(0);
	wire_y_pipeff_12_w_lg_w_q_range9344w9345w(0) <= NOT wire_y_pipeff_12_w_q_range9344w(0);
	wire_y_pipeff_12_w_lg_w_q_range9350w9351w(0) <= NOT wire_y_pipeff_12_w_q_range9350w(0);
	wire_y_pipeff_12_w_lg_w_q_range9356w9357w(0) <= NOT wire_y_pipeff_12_w_q_range9356w(0);
	wire_y_pipeff_12_w_lg_w_q_range9362w9363w(0) <= NOT wire_y_pipeff_12_w_q_range9362w(0);
	wire_y_pipeff_12_w_lg_w_q_range9368w9369w(0) <= NOT wire_y_pipeff_12_w_q_range9368w(0);
	wire_y_pipeff_12_w_lg_w_q_range9374w9375w(0) <= NOT wire_y_pipeff_12_w_q_range9374w(0);
	wire_y_pipeff_12_w_lg_w_q_range9380w9381w(0) <= NOT wire_y_pipeff_12_w_q_range9380w(0);
	wire_y_pipeff_12_w_lg_w_q_range9386w9387w(0) <= NOT wire_y_pipeff_12_w_q_range9386w(0);
	wire_y_pipeff_12_w_lg_w_q_range9392w9393w(0) <= NOT wire_y_pipeff_12_w_q_range9392w(0);
	wire_y_pipeff_12_w_lg_w_q_range9398w9399w(0) <= NOT wire_y_pipeff_12_w_q_range9398w(0);
	wire_y_pipeff_12_w_lg_w_q_range9404w9405w(0) <= NOT wire_y_pipeff_12_w_q_range9404w(0);
	wire_y_pipeff_12_w_lg_w_q_range9236w9237w(0) <= NOT wire_y_pipeff_12_w_q_range9236w(0);
	wire_y_pipeff_12_w_q_range9297w(0) <= y_pipeff_12(12);
	wire_y_pipeff_12_w_q_range9302w(0) <= y_pipeff_12(13);
	wire_y_pipeff_12_w_q_range9308w(0) <= y_pipeff_12(14);
	wire_y_pipeff_12_w_q_range9314w(0) <= y_pipeff_12(15);
	wire_y_pipeff_12_w_q_range9320w(0) <= y_pipeff_12(16);
	wire_y_pipeff_12_w_q_range9326w(0) <= y_pipeff_12(17);
	wire_y_pipeff_12_w_q_range9332w(0) <= y_pipeff_12(18);
	wire_y_pipeff_12_w_q_range9338w(0) <= y_pipeff_12(19);
	wire_y_pipeff_12_w_q_range9344w(0) <= y_pipeff_12(20);
	wire_y_pipeff_12_w_q_range9350w(0) <= y_pipeff_12(21);
	wire_y_pipeff_12_w_q_range9356w(0) <= y_pipeff_12(22);
	wire_y_pipeff_12_w_q_range9362w(0) <= y_pipeff_12(23);
	wire_y_pipeff_12_w_q_range9368w(0) <= y_pipeff_12(24);
	wire_y_pipeff_12_w_q_range9374w(0) <= y_pipeff_12(25);
	wire_y_pipeff_12_w_q_range9380w(0) <= y_pipeff_12(26);
	wire_y_pipeff_12_w_q_range9386w(0) <= y_pipeff_12(27);
	wire_y_pipeff_12_w_q_range9392w(0) <= y_pipeff_12(28);
	wire_y_pipeff_12_w_q_range9398w(0) <= y_pipeff_12(29);
	wire_y_pipeff_12_w_q_range9404w(0) <= y_pipeff_12(30);
	wire_y_pipeff_12_w_q_range9236w(0) <= y_pipeff_12(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_13 <= y_pipenode_13_w;
			END IF;
		END IF;
	END PROCESS;
	loop34 : FOR i IN 0 TO 31 GENERATE 
		wire_y_pipeff_13_w_lg_q9983w(i) <= y_pipeff_13(i) AND wire_sincosbitff_w_lg_w_q_range535w9982w(0);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 31 GENERATE 
		wire_y_pipeff_13_w_lg_q9986w(i) <= y_pipeff_13(i) AND wire_sincosbitff_w_q_range535w(0);
	END GENERATE loop35;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_2 <= y_pipenode_2_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_2_w_lg_w_q_range1569w1570w(0) <= NOT wire_y_pipeff_2_w_q_range1569w(0);
	wire_y_pipeff_2_w_lg_w_q_range1575w1576w(0) <= NOT wire_y_pipeff_2_w_q_range1575w(0);
	wire_y_pipeff_2_w_lg_w_q_range1581w1582w(0) <= NOT wire_y_pipeff_2_w_q_range1581w(0);
	wire_y_pipeff_2_w_lg_w_q_range1587w1588w(0) <= NOT wire_y_pipeff_2_w_q_range1587w(0);
	wire_y_pipeff_2_w_lg_w_q_range1593w1594w(0) <= NOT wire_y_pipeff_2_w_q_range1593w(0);
	wire_y_pipeff_2_w_lg_w_q_range1599w1600w(0) <= NOT wire_y_pipeff_2_w_q_range1599w(0);
	wire_y_pipeff_2_w_lg_w_q_range1605w1606w(0) <= NOT wire_y_pipeff_2_w_q_range1605w(0);
	wire_y_pipeff_2_w_lg_w_q_range1611w1612w(0) <= NOT wire_y_pipeff_2_w_q_range1611w(0);
	wire_y_pipeff_2_w_lg_w_q_range1617w1618w(0) <= NOT wire_y_pipeff_2_w_q_range1617w(0);
	wire_y_pipeff_2_w_lg_w_q_range1623w1624w(0) <= NOT wire_y_pipeff_2_w_q_range1623w(0);
	wire_y_pipeff_2_w_lg_w_q_range1629w1630w(0) <= NOT wire_y_pipeff_2_w_q_range1629w(0);
	wire_y_pipeff_2_w_lg_w_q_range1635w1636w(0) <= NOT wire_y_pipeff_2_w_q_range1635w(0);
	wire_y_pipeff_2_w_lg_w_q_range1641w1642w(0) <= NOT wire_y_pipeff_2_w_q_range1641w(0);
	wire_y_pipeff_2_w_lg_w_q_range1647w1648w(0) <= NOT wire_y_pipeff_2_w_q_range1647w(0);
	wire_y_pipeff_2_w_lg_w_q_range1653w1654w(0) <= NOT wire_y_pipeff_2_w_q_range1653w(0);
	wire_y_pipeff_2_w_lg_w_q_range1659w1660w(0) <= NOT wire_y_pipeff_2_w_q_range1659w(0);
	wire_y_pipeff_2_w_lg_w_q_range1665w1666w(0) <= NOT wire_y_pipeff_2_w_q_range1665w(0);
	wire_y_pipeff_2_w_lg_w_q_range1671w1672w(0) <= NOT wire_y_pipeff_2_w_q_range1671w(0);
	wire_y_pipeff_2_w_lg_w_q_range1677w1678w(0) <= NOT wire_y_pipeff_2_w_q_range1677w(0);
	wire_y_pipeff_2_w_lg_w_q_range1683w1684w(0) <= NOT wire_y_pipeff_2_w_q_range1683w(0);
	wire_y_pipeff_2_w_lg_w_q_range1522w1523w(0) <= NOT wire_y_pipeff_2_w_q_range1522w(0);
	wire_y_pipeff_2_w_lg_w_q_range1689w1690w(0) <= NOT wire_y_pipeff_2_w_q_range1689w(0);
	wire_y_pipeff_2_w_lg_w_q_range1501w1502w(0) <= NOT wire_y_pipeff_2_w_q_range1501w(0);
	wire_y_pipeff_2_w_lg_w_q_range1527w1528w(0) <= NOT wire_y_pipeff_2_w_q_range1527w(0);
	wire_y_pipeff_2_w_lg_w_q_range1533w1534w(0) <= NOT wire_y_pipeff_2_w_q_range1533w(0);
	wire_y_pipeff_2_w_lg_w_q_range1539w1540w(0) <= NOT wire_y_pipeff_2_w_q_range1539w(0);
	wire_y_pipeff_2_w_lg_w_q_range1545w1546w(0) <= NOT wire_y_pipeff_2_w_q_range1545w(0);
	wire_y_pipeff_2_w_lg_w_q_range1551w1552w(0) <= NOT wire_y_pipeff_2_w_q_range1551w(0);
	wire_y_pipeff_2_w_lg_w_q_range1557w1558w(0) <= NOT wire_y_pipeff_2_w_q_range1557w(0);
	wire_y_pipeff_2_w_lg_w_q_range1563w1564w(0) <= NOT wire_y_pipeff_2_w_q_range1563w(0);
	wire_y_pipeff_2_w_q_range1569w(0) <= y_pipeff_2(10);
	wire_y_pipeff_2_w_q_range1575w(0) <= y_pipeff_2(11);
	wire_y_pipeff_2_w_q_range1581w(0) <= y_pipeff_2(12);
	wire_y_pipeff_2_w_q_range1587w(0) <= y_pipeff_2(13);
	wire_y_pipeff_2_w_q_range1593w(0) <= y_pipeff_2(14);
	wire_y_pipeff_2_w_q_range1599w(0) <= y_pipeff_2(15);
	wire_y_pipeff_2_w_q_range1605w(0) <= y_pipeff_2(16);
	wire_y_pipeff_2_w_q_range1611w(0) <= y_pipeff_2(17);
	wire_y_pipeff_2_w_q_range1617w(0) <= y_pipeff_2(18);
	wire_y_pipeff_2_w_q_range1623w(0) <= y_pipeff_2(19);
	wire_y_pipeff_2_w_q_range1629w(0) <= y_pipeff_2(20);
	wire_y_pipeff_2_w_q_range1635w(0) <= y_pipeff_2(21);
	wire_y_pipeff_2_w_q_range1641w(0) <= y_pipeff_2(22);
	wire_y_pipeff_2_w_q_range1647w(0) <= y_pipeff_2(23);
	wire_y_pipeff_2_w_q_range1653w(0) <= y_pipeff_2(24);
	wire_y_pipeff_2_w_q_range1659w(0) <= y_pipeff_2(25);
	wire_y_pipeff_2_w_q_range1665w(0) <= y_pipeff_2(26);
	wire_y_pipeff_2_w_q_range1671w(0) <= y_pipeff_2(27);
	wire_y_pipeff_2_w_q_range1677w(0) <= y_pipeff_2(28);
	wire_y_pipeff_2_w_q_range1683w(0) <= y_pipeff_2(29);
	wire_y_pipeff_2_w_q_range1522w(0) <= y_pipeff_2(2);
	wire_y_pipeff_2_w_q_range1689w(0) <= y_pipeff_2(30);
	wire_y_pipeff_2_w_q_range1501w(0) <= y_pipeff_2(31);
	wire_y_pipeff_2_w_q_range1527w(0) <= y_pipeff_2(3);
	wire_y_pipeff_2_w_q_range1533w(0) <= y_pipeff_2(4);
	wire_y_pipeff_2_w_q_range1539w(0) <= y_pipeff_2(5);
	wire_y_pipeff_2_w_q_range1545w(0) <= y_pipeff_2(6);
	wire_y_pipeff_2_w_q_range1551w(0) <= y_pipeff_2(7);
	wire_y_pipeff_2_w_q_range1557w(0) <= y_pipeff_2(8);
	wire_y_pipeff_2_w_q_range1563w(0) <= y_pipeff_2(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_3 <= y_pipenode_3_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_3_w_lg_w_q_range2363w2364w(0) <= NOT wire_y_pipeff_3_w_q_range2363w(0);
	wire_y_pipeff_3_w_lg_w_q_range2369w2370w(0) <= NOT wire_y_pipeff_3_w_q_range2369w(0);
	wire_y_pipeff_3_w_lg_w_q_range2375w2376w(0) <= NOT wire_y_pipeff_3_w_q_range2375w(0);
	wire_y_pipeff_3_w_lg_w_q_range2381w2382w(0) <= NOT wire_y_pipeff_3_w_q_range2381w(0);
	wire_y_pipeff_3_w_lg_w_q_range2387w2388w(0) <= NOT wire_y_pipeff_3_w_q_range2387w(0);
	wire_y_pipeff_3_w_lg_w_q_range2393w2394w(0) <= NOT wire_y_pipeff_3_w_q_range2393w(0);
	wire_y_pipeff_3_w_lg_w_q_range2399w2400w(0) <= NOT wire_y_pipeff_3_w_q_range2399w(0);
	wire_y_pipeff_3_w_lg_w_q_range2405w2406w(0) <= NOT wire_y_pipeff_3_w_q_range2405w(0);
	wire_y_pipeff_3_w_lg_w_q_range2411w2412w(0) <= NOT wire_y_pipeff_3_w_q_range2411w(0);
	wire_y_pipeff_3_w_lg_w_q_range2417w2418w(0) <= NOT wire_y_pipeff_3_w_q_range2417w(0);
	wire_y_pipeff_3_w_lg_w_q_range2423w2424w(0) <= NOT wire_y_pipeff_3_w_q_range2423w(0);
	wire_y_pipeff_3_w_lg_w_q_range2429w2430w(0) <= NOT wire_y_pipeff_3_w_q_range2429w(0);
	wire_y_pipeff_3_w_lg_w_q_range2435w2436w(0) <= NOT wire_y_pipeff_3_w_q_range2435w(0);
	wire_y_pipeff_3_w_lg_w_q_range2441w2442w(0) <= NOT wire_y_pipeff_3_w_q_range2441w(0);
	wire_y_pipeff_3_w_lg_w_q_range2447w2448w(0) <= NOT wire_y_pipeff_3_w_q_range2447w(0);
	wire_y_pipeff_3_w_lg_w_q_range2453w2454w(0) <= NOT wire_y_pipeff_3_w_q_range2453w(0);
	wire_y_pipeff_3_w_lg_w_q_range2459w2460w(0) <= NOT wire_y_pipeff_3_w_q_range2459w(0);
	wire_y_pipeff_3_w_lg_w_q_range2465w2466w(0) <= NOT wire_y_pipeff_3_w_q_range2465w(0);
	wire_y_pipeff_3_w_lg_w_q_range2471w2472w(0) <= NOT wire_y_pipeff_3_w_q_range2471w(0);
	wire_y_pipeff_3_w_lg_w_q_range2477w2478w(0) <= NOT wire_y_pipeff_3_w_q_range2477w(0);
	wire_y_pipeff_3_w_lg_w_q_range2483w2484w(0) <= NOT wire_y_pipeff_3_w_q_range2483w(0);
	wire_y_pipeff_3_w_lg_w_q_range2297w2298w(0) <= NOT wire_y_pipeff_3_w_q_range2297w(0);
	wire_y_pipeff_3_w_lg_w_q_range2322w2323w(0) <= NOT wire_y_pipeff_3_w_q_range2322w(0);
	wire_y_pipeff_3_w_lg_w_q_range2327w2328w(0) <= NOT wire_y_pipeff_3_w_q_range2327w(0);
	wire_y_pipeff_3_w_lg_w_q_range2333w2334w(0) <= NOT wire_y_pipeff_3_w_q_range2333w(0);
	wire_y_pipeff_3_w_lg_w_q_range2339w2340w(0) <= NOT wire_y_pipeff_3_w_q_range2339w(0);
	wire_y_pipeff_3_w_lg_w_q_range2345w2346w(0) <= NOT wire_y_pipeff_3_w_q_range2345w(0);
	wire_y_pipeff_3_w_lg_w_q_range2351w2352w(0) <= NOT wire_y_pipeff_3_w_q_range2351w(0);
	wire_y_pipeff_3_w_lg_w_q_range2357w2358w(0) <= NOT wire_y_pipeff_3_w_q_range2357w(0);
	wire_y_pipeff_3_w_q_range2363w(0) <= y_pipeff_3(10);
	wire_y_pipeff_3_w_q_range2369w(0) <= y_pipeff_3(11);
	wire_y_pipeff_3_w_q_range2375w(0) <= y_pipeff_3(12);
	wire_y_pipeff_3_w_q_range2381w(0) <= y_pipeff_3(13);
	wire_y_pipeff_3_w_q_range2387w(0) <= y_pipeff_3(14);
	wire_y_pipeff_3_w_q_range2393w(0) <= y_pipeff_3(15);
	wire_y_pipeff_3_w_q_range2399w(0) <= y_pipeff_3(16);
	wire_y_pipeff_3_w_q_range2405w(0) <= y_pipeff_3(17);
	wire_y_pipeff_3_w_q_range2411w(0) <= y_pipeff_3(18);
	wire_y_pipeff_3_w_q_range2417w(0) <= y_pipeff_3(19);
	wire_y_pipeff_3_w_q_range2423w(0) <= y_pipeff_3(20);
	wire_y_pipeff_3_w_q_range2429w(0) <= y_pipeff_3(21);
	wire_y_pipeff_3_w_q_range2435w(0) <= y_pipeff_3(22);
	wire_y_pipeff_3_w_q_range2441w(0) <= y_pipeff_3(23);
	wire_y_pipeff_3_w_q_range2447w(0) <= y_pipeff_3(24);
	wire_y_pipeff_3_w_q_range2453w(0) <= y_pipeff_3(25);
	wire_y_pipeff_3_w_q_range2459w(0) <= y_pipeff_3(26);
	wire_y_pipeff_3_w_q_range2465w(0) <= y_pipeff_3(27);
	wire_y_pipeff_3_w_q_range2471w(0) <= y_pipeff_3(28);
	wire_y_pipeff_3_w_q_range2477w(0) <= y_pipeff_3(29);
	wire_y_pipeff_3_w_q_range2483w(0) <= y_pipeff_3(30);
	wire_y_pipeff_3_w_q_range2297w(0) <= y_pipeff_3(31);
	wire_y_pipeff_3_w_q_range2322w(0) <= y_pipeff_3(3);
	wire_y_pipeff_3_w_q_range2327w(0) <= y_pipeff_3(4);
	wire_y_pipeff_3_w_q_range2333w(0) <= y_pipeff_3(5);
	wire_y_pipeff_3_w_q_range2339w(0) <= y_pipeff_3(6);
	wire_y_pipeff_3_w_q_range2345w(0) <= y_pipeff_3(7);
	wire_y_pipeff_3_w_q_range2351w(0) <= y_pipeff_3(8);
	wire_y_pipeff_3_w_q_range2357w(0) <= y_pipeff_3(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_4 <= y_pipenode_4_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_4_w_lg_w_q_range3152w3153w(0) <= NOT wire_y_pipeff_4_w_q_range3152w(0);
	wire_y_pipeff_4_w_lg_w_q_range3158w3159w(0) <= NOT wire_y_pipeff_4_w_q_range3158w(0);
	wire_y_pipeff_4_w_lg_w_q_range3164w3165w(0) <= NOT wire_y_pipeff_4_w_q_range3164w(0);
	wire_y_pipeff_4_w_lg_w_q_range3170w3171w(0) <= NOT wire_y_pipeff_4_w_q_range3170w(0);
	wire_y_pipeff_4_w_lg_w_q_range3176w3177w(0) <= NOT wire_y_pipeff_4_w_q_range3176w(0);
	wire_y_pipeff_4_w_lg_w_q_range3182w3183w(0) <= NOT wire_y_pipeff_4_w_q_range3182w(0);
	wire_y_pipeff_4_w_lg_w_q_range3188w3189w(0) <= NOT wire_y_pipeff_4_w_q_range3188w(0);
	wire_y_pipeff_4_w_lg_w_q_range3194w3195w(0) <= NOT wire_y_pipeff_4_w_q_range3194w(0);
	wire_y_pipeff_4_w_lg_w_q_range3200w3201w(0) <= NOT wire_y_pipeff_4_w_q_range3200w(0);
	wire_y_pipeff_4_w_lg_w_q_range3206w3207w(0) <= NOT wire_y_pipeff_4_w_q_range3206w(0);
	wire_y_pipeff_4_w_lg_w_q_range3212w3213w(0) <= NOT wire_y_pipeff_4_w_q_range3212w(0);
	wire_y_pipeff_4_w_lg_w_q_range3218w3219w(0) <= NOT wire_y_pipeff_4_w_q_range3218w(0);
	wire_y_pipeff_4_w_lg_w_q_range3224w3225w(0) <= NOT wire_y_pipeff_4_w_q_range3224w(0);
	wire_y_pipeff_4_w_lg_w_q_range3230w3231w(0) <= NOT wire_y_pipeff_4_w_q_range3230w(0);
	wire_y_pipeff_4_w_lg_w_q_range3236w3237w(0) <= NOT wire_y_pipeff_4_w_q_range3236w(0);
	wire_y_pipeff_4_w_lg_w_q_range3242w3243w(0) <= NOT wire_y_pipeff_4_w_q_range3242w(0);
	wire_y_pipeff_4_w_lg_w_q_range3248w3249w(0) <= NOT wire_y_pipeff_4_w_q_range3248w(0);
	wire_y_pipeff_4_w_lg_w_q_range3254w3255w(0) <= NOT wire_y_pipeff_4_w_q_range3254w(0);
	wire_y_pipeff_4_w_lg_w_q_range3260w3261w(0) <= NOT wire_y_pipeff_4_w_q_range3260w(0);
	wire_y_pipeff_4_w_lg_w_q_range3266w3267w(0) <= NOT wire_y_pipeff_4_w_q_range3266w(0);
	wire_y_pipeff_4_w_lg_w_q_range3272w3273w(0) <= NOT wire_y_pipeff_4_w_q_range3272w(0);
	wire_y_pipeff_4_w_lg_w_q_range3088w3089w(0) <= NOT wire_y_pipeff_4_w_q_range3088w(0);
	wire_y_pipeff_4_w_lg_w_q_range3117w3118w(0) <= NOT wire_y_pipeff_4_w_q_range3117w(0);
	wire_y_pipeff_4_w_lg_w_q_range3122w3123w(0) <= NOT wire_y_pipeff_4_w_q_range3122w(0);
	wire_y_pipeff_4_w_lg_w_q_range3128w3129w(0) <= NOT wire_y_pipeff_4_w_q_range3128w(0);
	wire_y_pipeff_4_w_lg_w_q_range3134w3135w(0) <= NOT wire_y_pipeff_4_w_q_range3134w(0);
	wire_y_pipeff_4_w_lg_w_q_range3140w3141w(0) <= NOT wire_y_pipeff_4_w_q_range3140w(0);
	wire_y_pipeff_4_w_lg_w_q_range3146w3147w(0) <= NOT wire_y_pipeff_4_w_q_range3146w(0);
	wire_y_pipeff_4_w_q_range3152w(0) <= y_pipeff_4(10);
	wire_y_pipeff_4_w_q_range3158w(0) <= y_pipeff_4(11);
	wire_y_pipeff_4_w_q_range3164w(0) <= y_pipeff_4(12);
	wire_y_pipeff_4_w_q_range3170w(0) <= y_pipeff_4(13);
	wire_y_pipeff_4_w_q_range3176w(0) <= y_pipeff_4(14);
	wire_y_pipeff_4_w_q_range3182w(0) <= y_pipeff_4(15);
	wire_y_pipeff_4_w_q_range3188w(0) <= y_pipeff_4(16);
	wire_y_pipeff_4_w_q_range3194w(0) <= y_pipeff_4(17);
	wire_y_pipeff_4_w_q_range3200w(0) <= y_pipeff_4(18);
	wire_y_pipeff_4_w_q_range3206w(0) <= y_pipeff_4(19);
	wire_y_pipeff_4_w_q_range3212w(0) <= y_pipeff_4(20);
	wire_y_pipeff_4_w_q_range3218w(0) <= y_pipeff_4(21);
	wire_y_pipeff_4_w_q_range3224w(0) <= y_pipeff_4(22);
	wire_y_pipeff_4_w_q_range3230w(0) <= y_pipeff_4(23);
	wire_y_pipeff_4_w_q_range3236w(0) <= y_pipeff_4(24);
	wire_y_pipeff_4_w_q_range3242w(0) <= y_pipeff_4(25);
	wire_y_pipeff_4_w_q_range3248w(0) <= y_pipeff_4(26);
	wire_y_pipeff_4_w_q_range3254w(0) <= y_pipeff_4(27);
	wire_y_pipeff_4_w_q_range3260w(0) <= y_pipeff_4(28);
	wire_y_pipeff_4_w_q_range3266w(0) <= y_pipeff_4(29);
	wire_y_pipeff_4_w_q_range3272w(0) <= y_pipeff_4(30);
	wire_y_pipeff_4_w_q_range3088w(0) <= y_pipeff_4(31);
	wire_y_pipeff_4_w_q_range3117w(0) <= y_pipeff_4(4);
	wire_y_pipeff_4_w_q_range3122w(0) <= y_pipeff_4(5);
	wire_y_pipeff_4_w_q_range3128w(0) <= y_pipeff_4(6);
	wire_y_pipeff_4_w_q_range3134w(0) <= y_pipeff_4(7);
	wire_y_pipeff_4_w_q_range3140w(0) <= y_pipeff_4(8);
	wire_y_pipeff_4_w_q_range3146w(0) <= y_pipeff_4(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_5 <= y_pipenode_5_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_5_w_lg_w_q_range3936w3937w(0) <= NOT wire_y_pipeff_5_w_q_range3936w(0);
	wire_y_pipeff_5_w_lg_w_q_range3942w3943w(0) <= NOT wire_y_pipeff_5_w_q_range3942w(0);
	wire_y_pipeff_5_w_lg_w_q_range3948w3949w(0) <= NOT wire_y_pipeff_5_w_q_range3948w(0);
	wire_y_pipeff_5_w_lg_w_q_range3954w3955w(0) <= NOT wire_y_pipeff_5_w_q_range3954w(0);
	wire_y_pipeff_5_w_lg_w_q_range3960w3961w(0) <= NOT wire_y_pipeff_5_w_q_range3960w(0);
	wire_y_pipeff_5_w_lg_w_q_range3966w3967w(0) <= NOT wire_y_pipeff_5_w_q_range3966w(0);
	wire_y_pipeff_5_w_lg_w_q_range3972w3973w(0) <= NOT wire_y_pipeff_5_w_q_range3972w(0);
	wire_y_pipeff_5_w_lg_w_q_range3978w3979w(0) <= NOT wire_y_pipeff_5_w_q_range3978w(0);
	wire_y_pipeff_5_w_lg_w_q_range3984w3985w(0) <= NOT wire_y_pipeff_5_w_q_range3984w(0);
	wire_y_pipeff_5_w_lg_w_q_range3990w3991w(0) <= NOT wire_y_pipeff_5_w_q_range3990w(0);
	wire_y_pipeff_5_w_lg_w_q_range3996w3997w(0) <= NOT wire_y_pipeff_5_w_q_range3996w(0);
	wire_y_pipeff_5_w_lg_w_q_range4002w4003w(0) <= NOT wire_y_pipeff_5_w_q_range4002w(0);
	wire_y_pipeff_5_w_lg_w_q_range4008w4009w(0) <= NOT wire_y_pipeff_5_w_q_range4008w(0);
	wire_y_pipeff_5_w_lg_w_q_range4014w4015w(0) <= NOT wire_y_pipeff_5_w_q_range4014w(0);
	wire_y_pipeff_5_w_lg_w_q_range4020w4021w(0) <= NOT wire_y_pipeff_5_w_q_range4020w(0);
	wire_y_pipeff_5_w_lg_w_q_range4026w4027w(0) <= NOT wire_y_pipeff_5_w_q_range4026w(0);
	wire_y_pipeff_5_w_lg_w_q_range4032w4033w(0) <= NOT wire_y_pipeff_5_w_q_range4032w(0);
	wire_y_pipeff_5_w_lg_w_q_range4038w4039w(0) <= NOT wire_y_pipeff_5_w_q_range4038w(0);
	wire_y_pipeff_5_w_lg_w_q_range4044w4045w(0) <= NOT wire_y_pipeff_5_w_q_range4044w(0);
	wire_y_pipeff_5_w_lg_w_q_range4050w4051w(0) <= NOT wire_y_pipeff_5_w_q_range4050w(0);
	wire_y_pipeff_5_w_lg_w_q_range4056w4057w(0) <= NOT wire_y_pipeff_5_w_q_range4056w(0);
	wire_y_pipeff_5_w_lg_w_q_range3874w3875w(0) <= NOT wire_y_pipeff_5_w_q_range3874w(0);
	wire_y_pipeff_5_w_lg_w_q_range3907w3908w(0) <= NOT wire_y_pipeff_5_w_q_range3907w(0);
	wire_y_pipeff_5_w_lg_w_q_range3912w3913w(0) <= NOT wire_y_pipeff_5_w_q_range3912w(0);
	wire_y_pipeff_5_w_lg_w_q_range3918w3919w(0) <= NOT wire_y_pipeff_5_w_q_range3918w(0);
	wire_y_pipeff_5_w_lg_w_q_range3924w3925w(0) <= NOT wire_y_pipeff_5_w_q_range3924w(0);
	wire_y_pipeff_5_w_lg_w_q_range3930w3931w(0) <= NOT wire_y_pipeff_5_w_q_range3930w(0);
	wire_y_pipeff_5_w_q_range3936w(0) <= y_pipeff_5(10);
	wire_y_pipeff_5_w_q_range3942w(0) <= y_pipeff_5(11);
	wire_y_pipeff_5_w_q_range3948w(0) <= y_pipeff_5(12);
	wire_y_pipeff_5_w_q_range3954w(0) <= y_pipeff_5(13);
	wire_y_pipeff_5_w_q_range3960w(0) <= y_pipeff_5(14);
	wire_y_pipeff_5_w_q_range3966w(0) <= y_pipeff_5(15);
	wire_y_pipeff_5_w_q_range3972w(0) <= y_pipeff_5(16);
	wire_y_pipeff_5_w_q_range3978w(0) <= y_pipeff_5(17);
	wire_y_pipeff_5_w_q_range3984w(0) <= y_pipeff_5(18);
	wire_y_pipeff_5_w_q_range3990w(0) <= y_pipeff_5(19);
	wire_y_pipeff_5_w_q_range3996w(0) <= y_pipeff_5(20);
	wire_y_pipeff_5_w_q_range4002w(0) <= y_pipeff_5(21);
	wire_y_pipeff_5_w_q_range4008w(0) <= y_pipeff_5(22);
	wire_y_pipeff_5_w_q_range4014w(0) <= y_pipeff_5(23);
	wire_y_pipeff_5_w_q_range4020w(0) <= y_pipeff_5(24);
	wire_y_pipeff_5_w_q_range4026w(0) <= y_pipeff_5(25);
	wire_y_pipeff_5_w_q_range4032w(0) <= y_pipeff_5(26);
	wire_y_pipeff_5_w_q_range4038w(0) <= y_pipeff_5(27);
	wire_y_pipeff_5_w_q_range4044w(0) <= y_pipeff_5(28);
	wire_y_pipeff_5_w_q_range4050w(0) <= y_pipeff_5(29);
	wire_y_pipeff_5_w_q_range4056w(0) <= y_pipeff_5(30);
	wire_y_pipeff_5_w_q_range3874w(0) <= y_pipeff_5(31);
	wire_y_pipeff_5_w_q_range3907w(0) <= y_pipeff_5(5);
	wire_y_pipeff_5_w_q_range3912w(0) <= y_pipeff_5(6);
	wire_y_pipeff_5_w_q_range3918w(0) <= y_pipeff_5(7);
	wire_y_pipeff_5_w_q_range3924w(0) <= y_pipeff_5(8);
	wire_y_pipeff_5_w_q_range3930w(0) <= y_pipeff_5(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_6 <= y_pipenode_6_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_6_w_lg_w_q_range4715w4716w(0) <= NOT wire_y_pipeff_6_w_q_range4715w(0);
	wire_y_pipeff_6_w_lg_w_q_range4721w4722w(0) <= NOT wire_y_pipeff_6_w_q_range4721w(0);
	wire_y_pipeff_6_w_lg_w_q_range4727w4728w(0) <= NOT wire_y_pipeff_6_w_q_range4727w(0);
	wire_y_pipeff_6_w_lg_w_q_range4733w4734w(0) <= NOT wire_y_pipeff_6_w_q_range4733w(0);
	wire_y_pipeff_6_w_lg_w_q_range4739w4740w(0) <= NOT wire_y_pipeff_6_w_q_range4739w(0);
	wire_y_pipeff_6_w_lg_w_q_range4745w4746w(0) <= NOT wire_y_pipeff_6_w_q_range4745w(0);
	wire_y_pipeff_6_w_lg_w_q_range4751w4752w(0) <= NOT wire_y_pipeff_6_w_q_range4751w(0);
	wire_y_pipeff_6_w_lg_w_q_range4757w4758w(0) <= NOT wire_y_pipeff_6_w_q_range4757w(0);
	wire_y_pipeff_6_w_lg_w_q_range4763w4764w(0) <= NOT wire_y_pipeff_6_w_q_range4763w(0);
	wire_y_pipeff_6_w_lg_w_q_range4769w4770w(0) <= NOT wire_y_pipeff_6_w_q_range4769w(0);
	wire_y_pipeff_6_w_lg_w_q_range4775w4776w(0) <= NOT wire_y_pipeff_6_w_q_range4775w(0);
	wire_y_pipeff_6_w_lg_w_q_range4781w4782w(0) <= NOT wire_y_pipeff_6_w_q_range4781w(0);
	wire_y_pipeff_6_w_lg_w_q_range4787w4788w(0) <= NOT wire_y_pipeff_6_w_q_range4787w(0);
	wire_y_pipeff_6_w_lg_w_q_range4793w4794w(0) <= NOT wire_y_pipeff_6_w_q_range4793w(0);
	wire_y_pipeff_6_w_lg_w_q_range4799w4800w(0) <= NOT wire_y_pipeff_6_w_q_range4799w(0);
	wire_y_pipeff_6_w_lg_w_q_range4805w4806w(0) <= NOT wire_y_pipeff_6_w_q_range4805w(0);
	wire_y_pipeff_6_w_lg_w_q_range4811w4812w(0) <= NOT wire_y_pipeff_6_w_q_range4811w(0);
	wire_y_pipeff_6_w_lg_w_q_range4817w4818w(0) <= NOT wire_y_pipeff_6_w_q_range4817w(0);
	wire_y_pipeff_6_w_lg_w_q_range4823w4824w(0) <= NOT wire_y_pipeff_6_w_q_range4823w(0);
	wire_y_pipeff_6_w_lg_w_q_range4829w4830w(0) <= NOT wire_y_pipeff_6_w_q_range4829w(0);
	wire_y_pipeff_6_w_lg_w_q_range4835w4836w(0) <= NOT wire_y_pipeff_6_w_q_range4835w(0);
	wire_y_pipeff_6_w_lg_w_q_range4655w4656w(0) <= NOT wire_y_pipeff_6_w_q_range4655w(0);
	wire_y_pipeff_6_w_lg_w_q_range4692w4693w(0) <= NOT wire_y_pipeff_6_w_q_range4692w(0);
	wire_y_pipeff_6_w_lg_w_q_range4697w4698w(0) <= NOT wire_y_pipeff_6_w_q_range4697w(0);
	wire_y_pipeff_6_w_lg_w_q_range4703w4704w(0) <= NOT wire_y_pipeff_6_w_q_range4703w(0);
	wire_y_pipeff_6_w_lg_w_q_range4709w4710w(0) <= NOT wire_y_pipeff_6_w_q_range4709w(0);
	wire_y_pipeff_6_w_q_range4715w(0) <= y_pipeff_6(10);
	wire_y_pipeff_6_w_q_range4721w(0) <= y_pipeff_6(11);
	wire_y_pipeff_6_w_q_range4727w(0) <= y_pipeff_6(12);
	wire_y_pipeff_6_w_q_range4733w(0) <= y_pipeff_6(13);
	wire_y_pipeff_6_w_q_range4739w(0) <= y_pipeff_6(14);
	wire_y_pipeff_6_w_q_range4745w(0) <= y_pipeff_6(15);
	wire_y_pipeff_6_w_q_range4751w(0) <= y_pipeff_6(16);
	wire_y_pipeff_6_w_q_range4757w(0) <= y_pipeff_6(17);
	wire_y_pipeff_6_w_q_range4763w(0) <= y_pipeff_6(18);
	wire_y_pipeff_6_w_q_range4769w(0) <= y_pipeff_6(19);
	wire_y_pipeff_6_w_q_range4775w(0) <= y_pipeff_6(20);
	wire_y_pipeff_6_w_q_range4781w(0) <= y_pipeff_6(21);
	wire_y_pipeff_6_w_q_range4787w(0) <= y_pipeff_6(22);
	wire_y_pipeff_6_w_q_range4793w(0) <= y_pipeff_6(23);
	wire_y_pipeff_6_w_q_range4799w(0) <= y_pipeff_6(24);
	wire_y_pipeff_6_w_q_range4805w(0) <= y_pipeff_6(25);
	wire_y_pipeff_6_w_q_range4811w(0) <= y_pipeff_6(26);
	wire_y_pipeff_6_w_q_range4817w(0) <= y_pipeff_6(27);
	wire_y_pipeff_6_w_q_range4823w(0) <= y_pipeff_6(28);
	wire_y_pipeff_6_w_q_range4829w(0) <= y_pipeff_6(29);
	wire_y_pipeff_6_w_q_range4835w(0) <= y_pipeff_6(30);
	wire_y_pipeff_6_w_q_range4655w(0) <= y_pipeff_6(31);
	wire_y_pipeff_6_w_q_range4692w(0) <= y_pipeff_6(6);
	wire_y_pipeff_6_w_q_range4697w(0) <= y_pipeff_6(7);
	wire_y_pipeff_6_w_q_range4703w(0) <= y_pipeff_6(8);
	wire_y_pipeff_6_w_q_range4709w(0) <= y_pipeff_6(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_7 <= y_pipenode_7_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_7_w_lg_w_q_range5489w5490w(0) <= NOT wire_y_pipeff_7_w_q_range5489w(0);
	wire_y_pipeff_7_w_lg_w_q_range5495w5496w(0) <= NOT wire_y_pipeff_7_w_q_range5495w(0);
	wire_y_pipeff_7_w_lg_w_q_range5501w5502w(0) <= NOT wire_y_pipeff_7_w_q_range5501w(0);
	wire_y_pipeff_7_w_lg_w_q_range5507w5508w(0) <= NOT wire_y_pipeff_7_w_q_range5507w(0);
	wire_y_pipeff_7_w_lg_w_q_range5513w5514w(0) <= NOT wire_y_pipeff_7_w_q_range5513w(0);
	wire_y_pipeff_7_w_lg_w_q_range5519w5520w(0) <= NOT wire_y_pipeff_7_w_q_range5519w(0);
	wire_y_pipeff_7_w_lg_w_q_range5525w5526w(0) <= NOT wire_y_pipeff_7_w_q_range5525w(0);
	wire_y_pipeff_7_w_lg_w_q_range5531w5532w(0) <= NOT wire_y_pipeff_7_w_q_range5531w(0);
	wire_y_pipeff_7_w_lg_w_q_range5537w5538w(0) <= NOT wire_y_pipeff_7_w_q_range5537w(0);
	wire_y_pipeff_7_w_lg_w_q_range5543w5544w(0) <= NOT wire_y_pipeff_7_w_q_range5543w(0);
	wire_y_pipeff_7_w_lg_w_q_range5549w5550w(0) <= NOT wire_y_pipeff_7_w_q_range5549w(0);
	wire_y_pipeff_7_w_lg_w_q_range5555w5556w(0) <= NOT wire_y_pipeff_7_w_q_range5555w(0);
	wire_y_pipeff_7_w_lg_w_q_range5561w5562w(0) <= NOT wire_y_pipeff_7_w_q_range5561w(0);
	wire_y_pipeff_7_w_lg_w_q_range5567w5568w(0) <= NOT wire_y_pipeff_7_w_q_range5567w(0);
	wire_y_pipeff_7_w_lg_w_q_range5573w5574w(0) <= NOT wire_y_pipeff_7_w_q_range5573w(0);
	wire_y_pipeff_7_w_lg_w_q_range5579w5580w(0) <= NOT wire_y_pipeff_7_w_q_range5579w(0);
	wire_y_pipeff_7_w_lg_w_q_range5585w5586w(0) <= NOT wire_y_pipeff_7_w_q_range5585w(0);
	wire_y_pipeff_7_w_lg_w_q_range5591w5592w(0) <= NOT wire_y_pipeff_7_w_q_range5591w(0);
	wire_y_pipeff_7_w_lg_w_q_range5597w5598w(0) <= NOT wire_y_pipeff_7_w_q_range5597w(0);
	wire_y_pipeff_7_w_lg_w_q_range5603w5604w(0) <= NOT wire_y_pipeff_7_w_q_range5603w(0);
	wire_y_pipeff_7_w_lg_w_q_range5609w5610w(0) <= NOT wire_y_pipeff_7_w_q_range5609w(0);
	wire_y_pipeff_7_w_lg_w_q_range5431w5432w(0) <= NOT wire_y_pipeff_7_w_q_range5431w(0);
	wire_y_pipeff_7_w_lg_w_q_range5472w5473w(0) <= NOT wire_y_pipeff_7_w_q_range5472w(0);
	wire_y_pipeff_7_w_lg_w_q_range5477w5478w(0) <= NOT wire_y_pipeff_7_w_q_range5477w(0);
	wire_y_pipeff_7_w_lg_w_q_range5483w5484w(0) <= NOT wire_y_pipeff_7_w_q_range5483w(0);
	wire_y_pipeff_7_w_q_range5489w(0) <= y_pipeff_7(10);
	wire_y_pipeff_7_w_q_range5495w(0) <= y_pipeff_7(11);
	wire_y_pipeff_7_w_q_range5501w(0) <= y_pipeff_7(12);
	wire_y_pipeff_7_w_q_range5507w(0) <= y_pipeff_7(13);
	wire_y_pipeff_7_w_q_range5513w(0) <= y_pipeff_7(14);
	wire_y_pipeff_7_w_q_range5519w(0) <= y_pipeff_7(15);
	wire_y_pipeff_7_w_q_range5525w(0) <= y_pipeff_7(16);
	wire_y_pipeff_7_w_q_range5531w(0) <= y_pipeff_7(17);
	wire_y_pipeff_7_w_q_range5537w(0) <= y_pipeff_7(18);
	wire_y_pipeff_7_w_q_range5543w(0) <= y_pipeff_7(19);
	wire_y_pipeff_7_w_q_range5549w(0) <= y_pipeff_7(20);
	wire_y_pipeff_7_w_q_range5555w(0) <= y_pipeff_7(21);
	wire_y_pipeff_7_w_q_range5561w(0) <= y_pipeff_7(22);
	wire_y_pipeff_7_w_q_range5567w(0) <= y_pipeff_7(23);
	wire_y_pipeff_7_w_q_range5573w(0) <= y_pipeff_7(24);
	wire_y_pipeff_7_w_q_range5579w(0) <= y_pipeff_7(25);
	wire_y_pipeff_7_w_q_range5585w(0) <= y_pipeff_7(26);
	wire_y_pipeff_7_w_q_range5591w(0) <= y_pipeff_7(27);
	wire_y_pipeff_7_w_q_range5597w(0) <= y_pipeff_7(28);
	wire_y_pipeff_7_w_q_range5603w(0) <= y_pipeff_7(29);
	wire_y_pipeff_7_w_q_range5609w(0) <= y_pipeff_7(30);
	wire_y_pipeff_7_w_q_range5431w(0) <= y_pipeff_7(31);
	wire_y_pipeff_7_w_q_range5472w(0) <= y_pipeff_7(7);
	wire_y_pipeff_7_w_q_range5477w(0) <= y_pipeff_7(8);
	wire_y_pipeff_7_w_q_range5483w(0) <= y_pipeff_7(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_8 <= y_pipenode_8_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_8_w_lg_w_q_range6258w6259w(0) <= NOT wire_y_pipeff_8_w_q_range6258w(0);
	wire_y_pipeff_8_w_lg_w_q_range6264w6265w(0) <= NOT wire_y_pipeff_8_w_q_range6264w(0);
	wire_y_pipeff_8_w_lg_w_q_range6270w6271w(0) <= NOT wire_y_pipeff_8_w_q_range6270w(0);
	wire_y_pipeff_8_w_lg_w_q_range6276w6277w(0) <= NOT wire_y_pipeff_8_w_q_range6276w(0);
	wire_y_pipeff_8_w_lg_w_q_range6282w6283w(0) <= NOT wire_y_pipeff_8_w_q_range6282w(0);
	wire_y_pipeff_8_w_lg_w_q_range6288w6289w(0) <= NOT wire_y_pipeff_8_w_q_range6288w(0);
	wire_y_pipeff_8_w_lg_w_q_range6294w6295w(0) <= NOT wire_y_pipeff_8_w_q_range6294w(0);
	wire_y_pipeff_8_w_lg_w_q_range6300w6301w(0) <= NOT wire_y_pipeff_8_w_q_range6300w(0);
	wire_y_pipeff_8_w_lg_w_q_range6306w6307w(0) <= NOT wire_y_pipeff_8_w_q_range6306w(0);
	wire_y_pipeff_8_w_lg_w_q_range6312w6313w(0) <= NOT wire_y_pipeff_8_w_q_range6312w(0);
	wire_y_pipeff_8_w_lg_w_q_range6318w6319w(0) <= NOT wire_y_pipeff_8_w_q_range6318w(0);
	wire_y_pipeff_8_w_lg_w_q_range6324w6325w(0) <= NOT wire_y_pipeff_8_w_q_range6324w(0);
	wire_y_pipeff_8_w_lg_w_q_range6330w6331w(0) <= NOT wire_y_pipeff_8_w_q_range6330w(0);
	wire_y_pipeff_8_w_lg_w_q_range6336w6337w(0) <= NOT wire_y_pipeff_8_w_q_range6336w(0);
	wire_y_pipeff_8_w_lg_w_q_range6342w6343w(0) <= NOT wire_y_pipeff_8_w_q_range6342w(0);
	wire_y_pipeff_8_w_lg_w_q_range6348w6349w(0) <= NOT wire_y_pipeff_8_w_q_range6348w(0);
	wire_y_pipeff_8_w_lg_w_q_range6354w6355w(0) <= NOT wire_y_pipeff_8_w_q_range6354w(0);
	wire_y_pipeff_8_w_lg_w_q_range6360w6361w(0) <= NOT wire_y_pipeff_8_w_q_range6360w(0);
	wire_y_pipeff_8_w_lg_w_q_range6366w6367w(0) <= NOT wire_y_pipeff_8_w_q_range6366w(0);
	wire_y_pipeff_8_w_lg_w_q_range6372w6373w(0) <= NOT wire_y_pipeff_8_w_q_range6372w(0);
	wire_y_pipeff_8_w_lg_w_q_range6378w6379w(0) <= NOT wire_y_pipeff_8_w_q_range6378w(0);
	wire_y_pipeff_8_w_lg_w_q_range6202w6203w(0) <= NOT wire_y_pipeff_8_w_q_range6202w(0);
	wire_y_pipeff_8_w_lg_w_q_range6247w6248w(0) <= NOT wire_y_pipeff_8_w_q_range6247w(0);
	wire_y_pipeff_8_w_lg_w_q_range6252w6253w(0) <= NOT wire_y_pipeff_8_w_q_range6252w(0);
	wire_y_pipeff_8_w_q_range6258w(0) <= y_pipeff_8(10);
	wire_y_pipeff_8_w_q_range6264w(0) <= y_pipeff_8(11);
	wire_y_pipeff_8_w_q_range6270w(0) <= y_pipeff_8(12);
	wire_y_pipeff_8_w_q_range6276w(0) <= y_pipeff_8(13);
	wire_y_pipeff_8_w_q_range6282w(0) <= y_pipeff_8(14);
	wire_y_pipeff_8_w_q_range6288w(0) <= y_pipeff_8(15);
	wire_y_pipeff_8_w_q_range6294w(0) <= y_pipeff_8(16);
	wire_y_pipeff_8_w_q_range6300w(0) <= y_pipeff_8(17);
	wire_y_pipeff_8_w_q_range6306w(0) <= y_pipeff_8(18);
	wire_y_pipeff_8_w_q_range6312w(0) <= y_pipeff_8(19);
	wire_y_pipeff_8_w_q_range6318w(0) <= y_pipeff_8(20);
	wire_y_pipeff_8_w_q_range6324w(0) <= y_pipeff_8(21);
	wire_y_pipeff_8_w_q_range6330w(0) <= y_pipeff_8(22);
	wire_y_pipeff_8_w_q_range6336w(0) <= y_pipeff_8(23);
	wire_y_pipeff_8_w_q_range6342w(0) <= y_pipeff_8(24);
	wire_y_pipeff_8_w_q_range6348w(0) <= y_pipeff_8(25);
	wire_y_pipeff_8_w_q_range6354w(0) <= y_pipeff_8(26);
	wire_y_pipeff_8_w_q_range6360w(0) <= y_pipeff_8(27);
	wire_y_pipeff_8_w_q_range6366w(0) <= y_pipeff_8(28);
	wire_y_pipeff_8_w_q_range6372w(0) <= y_pipeff_8(29);
	wire_y_pipeff_8_w_q_range6378w(0) <= y_pipeff_8(30);
	wire_y_pipeff_8_w_q_range6202w(0) <= y_pipeff_8(31);
	wire_y_pipeff_8_w_q_range6247w(0) <= y_pipeff_8(8);
	wire_y_pipeff_8_w_q_range6252w(0) <= y_pipeff_8(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN y_pipeff_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN y_pipeff_9 <= y_pipenode_9_w;
			END IF;
		END IF;
	END PROCESS;
	wire_y_pipeff_9_w_lg_w_q_range7022w7023w(0) <= NOT wire_y_pipeff_9_w_q_range7022w(0);
	wire_y_pipeff_9_w_lg_w_q_range7028w7029w(0) <= NOT wire_y_pipeff_9_w_q_range7028w(0);
	wire_y_pipeff_9_w_lg_w_q_range7034w7035w(0) <= NOT wire_y_pipeff_9_w_q_range7034w(0);
	wire_y_pipeff_9_w_lg_w_q_range7040w7041w(0) <= NOT wire_y_pipeff_9_w_q_range7040w(0);
	wire_y_pipeff_9_w_lg_w_q_range7046w7047w(0) <= NOT wire_y_pipeff_9_w_q_range7046w(0);
	wire_y_pipeff_9_w_lg_w_q_range7052w7053w(0) <= NOT wire_y_pipeff_9_w_q_range7052w(0);
	wire_y_pipeff_9_w_lg_w_q_range7058w7059w(0) <= NOT wire_y_pipeff_9_w_q_range7058w(0);
	wire_y_pipeff_9_w_lg_w_q_range7064w7065w(0) <= NOT wire_y_pipeff_9_w_q_range7064w(0);
	wire_y_pipeff_9_w_lg_w_q_range7070w7071w(0) <= NOT wire_y_pipeff_9_w_q_range7070w(0);
	wire_y_pipeff_9_w_lg_w_q_range7076w7077w(0) <= NOT wire_y_pipeff_9_w_q_range7076w(0);
	wire_y_pipeff_9_w_lg_w_q_range7082w7083w(0) <= NOT wire_y_pipeff_9_w_q_range7082w(0);
	wire_y_pipeff_9_w_lg_w_q_range7088w7089w(0) <= NOT wire_y_pipeff_9_w_q_range7088w(0);
	wire_y_pipeff_9_w_lg_w_q_range7094w7095w(0) <= NOT wire_y_pipeff_9_w_q_range7094w(0);
	wire_y_pipeff_9_w_lg_w_q_range7100w7101w(0) <= NOT wire_y_pipeff_9_w_q_range7100w(0);
	wire_y_pipeff_9_w_lg_w_q_range7106w7107w(0) <= NOT wire_y_pipeff_9_w_q_range7106w(0);
	wire_y_pipeff_9_w_lg_w_q_range7112w7113w(0) <= NOT wire_y_pipeff_9_w_q_range7112w(0);
	wire_y_pipeff_9_w_lg_w_q_range7118w7119w(0) <= NOT wire_y_pipeff_9_w_q_range7118w(0);
	wire_y_pipeff_9_w_lg_w_q_range7124w7125w(0) <= NOT wire_y_pipeff_9_w_q_range7124w(0);
	wire_y_pipeff_9_w_lg_w_q_range7130w7131w(0) <= NOT wire_y_pipeff_9_w_q_range7130w(0);
	wire_y_pipeff_9_w_lg_w_q_range7136w7137w(0) <= NOT wire_y_pipeff_9_w_q_range7136w(0);
	wire_y_pipeff_9_w_lg_w_q_range7142w7143w(0) <= NOT wire_y_pipeff_9_w_q_range7142w(0);
	wire_y_pipeff_9_w_lg_w_q_range6968w6969w(0) <= NOT wire_y_pipeff_9_w_q_range6968w(0);
	wire_y_pipeff_9_w_lg_w_q_range7017w7018w(0) <= NOT wire_y_pipeff_9_w_q_range7017w(0);
	wire_y_pipeff_9_w_q_range7022w(0) <= y_pipeff_9(10);
	wire_y_pipeff_9_w_q_range7028w(0) <= y_pipeff_9(11);
	wire_y_pipeff_9_w_q_range7034w(0) <= y_pipeff_9(12);
	wire_y_pipeff_9_w_q_range7040w(0) <= y_pipeff_9(13);
	wire_y_pipeff_9_w_q_range7046w(0) <= y_pipeff_9(14);
	wire_y_pipeff_9_w_q_range7052w(0) <= y_pipeff_9(15);
	wire_y_pipeff_9_w_q_range7058w(0) <= y_pipeff_9(16);
	wire_y_pipeff_9_w_q_range7064w(0) <= y_pipeff_9(17);
	wire_y_pipeff_9_w_q_range7070w(0) <= y_pipeff_9(18);
	wire_y_pipeff_9_w_q_range7076w(0) <= y_pipeff_9(19);
	wire_y_pipeff_9_w_q_range7082w(0) <= y_pipeff_9(20);
	wire_y_pipeff_9_w_q_range7088w(0) <= y_pipeff_9(21);
	wire_y_pipeff_9_w_q_range7094w(0) <= y_pipeff_9(22);
	wire_y_pipeff_9_w_q_range7100w(0) <= y_pipeff_9(23);
	wire_y_pipeff_9_w_q_range7106w(0) <= y_pipeff_9(24);
	wire_y_pipeff_9_w_q_range7112w(0) <= y_pipeff_9(25);
	wire_y_pipeff_9_w_q_range7118w(0) <= y_pipeff_9(26);
	wire_y_pipeff_9_w_q_range7124w(0) <= y_pipeff_9(27);
	wire_y_pipeff_9_w_q_range7130w(0) <= y_pipeff_9(28);
	wire_y_pipeff_9_w_q_range7136w(0) <= y_pipeff_9(29);
	wire_y_pipeff_9_w_q_range7142w(0) <= y_pipeff_9(30);
	wire_y_pipeff_9_w_q_range6968w(0) <= y_pipeff_9(31);
	wire_y_pipeff_9_w_q_range7017w(0) <= y_pipeff_9(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_0 <= radians_load_node_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_1 <= wire_z_pipeff1_sub_result;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_1_w_q_range1241w(0) <= z_pipeff_1(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_10 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_10 <= z_pipenode_10_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_10_w_q_range8225w(0) <= z_pipeff_10(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_11 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_11 <= z_pipenode_11_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_11_w_q_range8976w(0) <= z_pipeff_11(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_12 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_12 <= z_pipenode_12_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_12_w_q_range9722w(0) <= z_pipeff_12(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_13 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_13 <= z_pipenode_13_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_2 <= z_pipenode_2_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_2_w_q_range2037w(0) <= z_pipeff_2(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_3 <= z_pipenode_3_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_3_w_q_range2828w(0) <= z_pipeff_3(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_4 <= z_pipenode_4_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_4_w_q_range3614w(0) <= z_pipeff_4(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_5 <= z_pipenode_5_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_5_w_q_range4395w(0) <= z_pipeff_5(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_6 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_6 <= z_pipenode_6_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_6_w_q_range5171w(0) <= z_pipeff_6(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_7 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_7 <= z_pipenode_7_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_7_w_q_range5942w(0) <= z_pipeff_7(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_8 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_8 <= z_pipenode_8_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_8_w_q_range6708w(0) <= z_pipeff_8(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN z_pipeff_9 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN z_pipeff_9 <= z_pipenode_9_w;
			END IF;
		END IF;
	END PROCESS;
	wire_z_pipeff_9_w_q_range7469w(0) <= z_pipeff_9(31);
	wire_sincos_add_cin <= wire_sincosbitff_w_lg_w_q_range9989w9990w(0);
	sincos_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => wire_sincos_add_cin,
		dataa => delay_pipe_w,
		datab => post_estimate_w,
		result => wire_sincos_add_result
	  );
	x_pipenode_10_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_9(31),
		dataa => x_pipeff_9,
		datab => x_subnode_10_w,
		result => wire_x_pipenode_10_add_result
	  );
	x_pipenode_11_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_10(31),
		dataa => x_pipeff_10,
		datab => x_subnode_11_w,
		result => wire_x_pipenode_11_add_result
	  );
	x_pipenode_12_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_11(31),
		dataa => x_pipeff_11,
		datab => x_subnode_12_w,
		result => wire_x_pipenode_12_add_result
	  );
	x_pipenode_13_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_12(31),
		dataa => x_pipeff_12,
		datab => x_subnode_13_w,
		result => wire_x_pipenode_13_add_result
	  );
	x_pipenode_2_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_1(31),
		dataa => x_pipeff_1,
		datab => x_subnode_2_w,
		result => wire_x_pipenode_2_add_result
	  );
	x_pipenode_3_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_2(31),
		dataa => x_pipeff_2,
		datab => x_subnode_3_w,
		result => wire_x_pipenode_3_add_result
	  );
	x_pipenode_4_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_3(31),
		dataa => x_pipeff_3,
		datab => x_subnode_4_w,
		result => wire_x_pipenode_4_add_result
	  );
	x_pipenode_5_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_4(31),
		dataa => x_pipeff_4,
		datab => x_subnode_5_w,
		result => wire_x_pipenode_5_add_result
	  );
	x_pipenode_6_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_5(31),
		dataa => x_pipeff_5,
		datab => x_subnode_6_w,
		result => wire_x_pipenode_6_add_result
	  );
	x_pipenode_7_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_6(31),
		dataa => x_pipeff_6,
		datab => x_subnode_7_w,
		result => wire_x_pipenode_7_add_result
	  );
	x_pipenode_8_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_7(31),
		dataa => x_pipeff_7,
		datab => x_subnode_8_w,
		result => wire_x_pipenode_8_add_result
	  );
	x_pipenode_9_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_8(31),
		dataa => x_pipeff_8,
		datab => x_subnode_9_w,
		result => wire_x_pipenode_9_add_result
	  );
	y_pipeff1_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		dataa => y_pipeff_0,
		datab => y_subnode_1_w,
		result => wire_y_pipeff1_add_result
	  );
	y_pipenode_10_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_9(31),
		dataa => y_pipeff_9,
		datab => y_subnode_10_w,
		result => wire_y_pipenode_10_add_result
	  );
	y_pipenode_11_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_10(31),
		dataa => y_pipeff_10,
		datab => y_subnode_11_w,
		result => wire_y_pipenode_11_add_result
	  );
	y_pipenode_12_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_11(31),
		dataa => y_pipeff_11,
		datab => y_subnode_12_w,
		result => wire_y_pipenode_12_add_result
	  );
	y_pipenode_13_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_12(31),
		dataa => y_pipeff_12,
		datab => y_subnode_13_w,
		result => wire_y_pipenode_13_add_result
	  );
	y_pipenode_2_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_1(31),
		dataa => y_pipeff_1,
		datab => y_subnode_2_w,
		result => wire_y_pipenode_2_add_result
	  );
	y_pipenode_3_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_2(31),
		dataa => y_pipeff_2,
		datab => y_subnode_3_w,
		result => wire_y_pipenode_3_add_result
	  );
	y_pipenode_4_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_3(31),
		dataa => y_pipeff_3,
		datab => y_subnode_4_w,
		result => wire_y_pipenode_4_add_result
	  );
	y_pipenode_5_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_4(31),
		dataa => y_pipeff_4,
		datab => y_subnode_5_w,
		result => wire_y_pipenode_5_add_result
	  );
	y_pipenode_6_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_5(31),
		dataa => y_pipeff_5,
		datab => y_subnode_6_w,
		result => wire_y_pipenode_6_add_result
	  );
	y_pipenode_7_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_6(31),
		dataa => y_pipeff_6,
		datab => y_subnode_7_w,
		result => wire_y_pipenode_7_add_result
	  );
	y_pipenode_8_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_7(31),
		dataa => y_pipeff_7,
		datab => y_subnode_8_w,
		result => wire_y_pipenode_8_add_result
	  );
	y_pipenode_9_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_8(31),
		dataa => y_pipeff_8,
		datab => y_subnode_9_w,
		result => wire_y_pipenode_9_add_result
	  );
	z_pipeff1_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		dataa => z_pipeff_0,
		datab => atannode_0_w,
		result => wire_z_pipeff1_sub_result
	  );
	z_pipenode_10_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_9(31),
		dataa => z_pipeff_9,
		datab => z_subnode_10_w,
		result => wire_z_pipenode_10_add_result
	  );
	z_pipenode_11_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_10(31),
		dataa => z_pipeff_10,
		datab => z_subnode_11_w,
		result => wire_z_pipenode_11_add_result
	  );
	z_pipenode_12_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_11(31),
		dataa => z_pipeff_11,
		datab => z_subnode_12_w,
		result => wire_z_pipenode_12_add_result
	  );
	z_pipenode_13_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_12(31),
		dataa => z_pipeff_12,
		datab => z_subnode_13_w,
		result => wire_z_pipenode_13_add_result
	  );
	z_pipenode_2_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_1(31),
		dataa => z_pipeff_1,
		datab => z_subnode_2_w,
		result => wire_z_pipenode_2_add_result
	  );
	z_pipenode_3_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_2(31),
		dataa => z_pipeff_2,
		datab => z_subnode_3_w,
		result => wire_z_pipenode_3_add_result
	  );
	z_pipenode_4_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_3(31),
		dataa => z_pipeff_3,
		datab => z_subnode_4_w,
		result => wire_z_pipenode_4_add_result
	  );
	z_pipenode_5_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_4(31),
		dataa => z_pipeff_4,
		datab => z_subnode_5_w,
		result => wire_z_pipenode_5_add_result
	  );
	z_pipenode_6_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_5(31),
		dataa => z_pipeff_5,
		datab => z_subnode_6_w,
		result => wire_z_pipenode_6_add_result
	  );
	z_pipenode_7_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_6(31),
		dataa => z_pipeff_6,
		datab => z_subnode_7_w,
		result => wire_z_pipenode_7_add_result
	  );
	z_pipenode_8_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_7(31),
		dataa => z_pipeff_7,
		datab => z_subnode_8_w,
		result => wire_z_pipenode_8_add_result
	  );
	z_pipenode_9_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		cin => z_pipeff_8(31),
		dataa => z_pipeff_8,
		datab => z_subnode_9_w,
		result => wire_z_pipenode_9_add_result
	  );
	cmx :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTHA => 32,
		LPM_WIDTHB => 32,
		LPM_WIDTHP => 64
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => multiplier_input_w,
		datab => z_pipeff_13,
		result => wire_cmx_result
	  );

 END RTL; --coshw_altfp_sincos_cordic_m_d5e


--altfp_sincos_range CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" WIDTH_EXP=8 WIDTH_MAN=23 aclr circle clken clock data negcircle
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END


--altfp_sincos_srrt CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone V" address basefraction incexponent incmantissa
--VERSION_BEGIN 18.1 cbx_altfp_sincos 2018:09:12:13:04:24:SJ cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_cycloneii 2018:09:12:13:04:24:SJ cbx_lpm_add_sub 2018:09:12:13:04:24:SJ cbx_lpm_clshift 2018:09:12:13:04:24:SJ cbx_lpm_mult 2018:09:12:13:04:24:SJ cbx_lpm_mux 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ cbx_nadder 2018:09:12:13:04:24:SJ cbx_padd 2018:09:12:13:04:24:SJ cbx_stratix 2018:09:12:13:04:24:SJ cbx_stratixii 2018:09:12:13:04:24:SJ cbx_util_mgl 2018:09:12:13:04:24:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_mux 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_srrt_koa IS 
	 PORT 
	 ( 
		 address	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 basefraction	:	OUT  STD_LOGIC_VECTOR (35 DOWNTO 0);
		 incexponent	:	OUT  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 incmantissa	:	OUT  STD_LOGIC_VECTOR (55 DOWNTO 0)
	 ); 
 END coshw_altfp_sincos_srrt_koa;

 ARCHITECTURE RTL OF coshw_altfp_sincos_srrt_koa IS

	 SIGNAL  wire_mux2_data	:	STD_LOGIC_VECTOR (25599 DOWNTO 0);
	 SIGNAL  wire_mux2_data_2d	:	STD_LOGIC_2D(255 DOWNTO 0, 99 DOWNTO 0);
	 SIGNAL  wire_mux2_result	:	STD_LOGIC_VECTOR (99 DOWNTO 0);
 BEGIN

	basefraction <= wire_mux2_result(35 DOWNTO 0);
	incexponent <= wire_mux2_result(99 DOWNTO 92);
	incmantissa <= wire_mux2_result(91 DOWNTO 36);
	wire_mux2_data <= ( "00000000" & "10011010011011101110000001101101101100010100101011001000" & "00110110" & "1101100010100101011001100101" & "00000001" & "10011010011011101110000001101101101100010100101011010000" & "00011011" & "0110110001010010101100110010" & "00000000" & "10100110100110111011100000011011011011000101001010111000" & "00001101" & "1011011000101001010110011001" & "00000001" & "10100110100110111011100000011011011011000101001010110000" & "00000110" & "1101101100010100101011001101" & "00000000" & "10101001101001101110111000000110110110110001010010110000" & "00000011" & "0110110110001010010101100110" & "00000000" & "11010100110100110111011100000011011011011000101001100000" & "10000001" & "1011011011000101001010110011" & "00000000" & "11101010011010011011101110000001101101101100010100011000" & "11000000" & "1101101101100010100101011010" & "00000000" & "11110101001101001101110111000000110110110110001010011000" & "11100000" & "0110110110110001010010101101" & "00000000" & "11111010100110100110111011100000011011011011000101010000" & "01110000" & "0011011011011000101001010110" & "00000001" & "11111010100110100110111011100000011011011011000101010000" & "10111000" & "0001101101101100010100101011" & "00000010" & "11111010100110100110111011100000011011011011000101010000" & "11011100" & "0000110110110110001010010110" & "00000011" & "11111010100110100110111011100000011011011011000100101000" & "11101110" & "0000011011011011000101001011" & "00000000" & "10001111101010011010011011101110000001101101101100011000" & "01110111" & "0000001101101101100010100101" & "00000001" & "10001111101010011010011011101110000001101101101100100000" & "10111011" & "1000000110110110110001010011" & "00000000" & "10100011111010100110100110111011100000011011011011001000" & "11011101" & "1100000011011011011000101001" & "00000000" & "11010001111101010011010011011101110000001101101101010000" & "01101110" & "1110000001101101101100010101" & "00000000" & "11101000111110101001101001101110111000000110110110111000" & "00110111" & "0111000000110110110110001010"
 & "00000000" & "11110100011111010100110100110111011100000011011011011000" & "10011011" & "1011100000011011011011000101" & "00000000" & "11111010001111101010011010011011101110000001101101101000" & "01001101" & "1101110000001101101101100011" & "00000001" & "11111010001111101010011010011011101110000001101110000000" & "10100110" & "1110111000000110110110110001" & "00000000" & "10111110100011111010100110100110111011100000011011100000" & "11010011" & "0111011100000011011011011001" & "00000001" & "10111110100011111010100110100110111011100000011011101000" & "01101001" & "1011101110000001101101101100" & "00000000" & "10101111101000111110101001101001101110111000000110111000" & "00110100" & "1101110111000000110110110110" & "00000001" & "10101111101000111110101001101001101110111000000110110000" & "10011010" & "0110111011100000011011011011" & "00000000" & "10101011111010001111101010011010011011101110000001110000" & "01001101" & "0011011101110000001101101110" & "00000000" & "11010101111101000111110101001101001101110111000000111000" & "10100110" & "1001101110111000000110110111" & "00000000" & "11101010111110100011111010100110100110111011100000110000" & "01010011" & "0100110111011100000011011011" & "00000001" & "11101010111110100011111010100110100110111011100000100000" & "10101001" & "1010011011101110000001101110" & "00000010" & "11101010111110100011111010100110100110111011011111111000" & "11010100" & "1101001101110111000000110111" & "00000000" & "10011101010111110100011111010100110100110111011100000000" & "11101010" & "0110100110111011100000011011" & "00000001" & "10011101010111110100011111010100110100110111011100011000" & "11110101" & "0011010011011101110000001110" & "00000010" & "10011101010111110100011111010100110100110111011100011000" & "11111010" & "1001101001101110111000000111" & "00000011" & "10011101010111110100011111010100110100110111011100011000" & "01111101" & "0100110100110111011100000011" & "00000100" & "10011101010111110100011111010100110100110111011110010000" & "00111110" & "1010011010011011101110000010" & "00000000"
 & "10000100111010101111101000111110101001101001101111000000" & "00011111" & "0101001101001101110111000001" & "00000000" & "11000010011101010111110100011111010100110100110111011000" & "10001111" & "1010100110100110111011100000" & "00000000" & "11100001001110101011111010001111101010011010011011110000" & "01000111" & "1101010011010011011101110000" & "00000000" & "11110000100111010101111101000111110101001101001110000000" & "10100011" & "1110101001101001101110111000" & "00000000" & "11111000010011101010111110100011111010100110100110111000" & "11010001" & "1111010100110100110111011100" & "00000000" & "11111100001001110101011111010001111101010011010011011000" & "11101000" & "1111101010011010011011101110" & "00000000" & "11111110000100111010101111101000111110101001101001110000" & "11110100" & "0111110101001101001101110111" & "00000001" & "11111110000100111010101111101000111110101001101010000000" & "11111010" & "0011111010100110100110111100" & "00000010" & "11111110000100111010101111101000111110101001101001110000" & "01111101" & "0001111101010011010011011110" & "00000000" & "10011111110000100111010101111101000111110101001101011000" & "10111110" & "1000111110101001101001101111" & "00000001" & "10011111110000100111010101111101000111110101001101100000" & "01011111" & "0100011111010100110100110111" & "00000000" & "10100111111100001001110101011111010001111101010011010000" & "10101111" & "1010001111101010011010011100" & "00000001" & "10100111111100001001110101011111010001111101010011100000" & "01010111" & "1101000111110101001101001110" & "00000010" & "10100111111100001001110101011111010001111101010011010000" & "10101011" & "1110100011111010100110100111" & "00000000" & "10010100111111100001001110101011111010001111101010011000" & "11010101" & "1111010001111101010011010011" & "00000001" & "10010100111111100001001110101011111010001111101010101000" & "11101010" & "1111101000111110101001101010" & "00000000" & "10100101001111111000010011101010111110100011111010101000" & "01110101" & "0111110100011111010100110101" & "00000001" & "10100101001111111000010011101010111110100011111010101000"
 & "00111010" & "1011111010001111101010011010" & "00000000" & "10101001010011111110000100111010101111101000111110101000" & "10011101" & "0101111101000111110101001101" & "00000001" & "10101001010011111110000100111010101111101000111110111000" & "01001110" & "1010111110100011111010100111" & "00000010" & "10101001010011111110000100111010101111101000111110111000" & "00100111" & "0101011111010001111101010011" & "00000011" & "10101001010011111110000100111010101111101000111110111000" & "00010011" & "1010101111101000111110101010" & "00000100" & "10101001010011111110000100111010101111101000111110111000" & "00001001" & "1101010111110100011111010101" & "00000101" & "10101001010011111110000100111010101111101001000000110000" & "10000100" & "1110101011111010001111101010" & "00000000" & "10000010101001010011111110000100111010101111101001001000" & "11000010" & "0111010101111101000111110101" & "00000001" & "10000010101001010011111110000100111010101111101001010000" & "11100001" & "0011101010111110100011111011" & "00000010" & "10000010101001010011111110000100111010101111101000111000" & "11110000" & "1001110101011111010001111101" & "00000011" & "10000010101001010011111110000100111010101111101001100000" & "11111000" & "0100111010101111101000111111" & "00000000" & "10001000001010100101001111111000010011101010111110100000" & "11111100" & "0010011101010111110100011111" & "00000001" & "10001000001010100101001111111000010011101010111110100000" & "11111110" & "0001001110101011111010010000" & "00000010" & "10001000001010100101001111111000010011101010111110100000" & "01111111" & "0000100111010101111101001000" & "00000000" & "10010001000001010100101001111111000010011101011000010000" & "00111111" & "1000010011101010111110100100" & "00000000" & "11001000100000101010010100111111100001001110101011111000" & "10011111" & "1100001001110101011111010010" & "00000000" & "11100100010000010101001010011111110000100111010101111000" & "01001111" & "1110000100111010101111101001" & "00000001" & "11100100010000010101001010011111110000100111010101110000" & "10100111"
 & "1111000010011101010111110100" & "00000010" & "11100100010000010101001010011111110000100111010110001000" & "01010011" & "1111100001001110101011111010" & "00000000" & "10011100100010000010101001010011111110000100111010111000" & "00101001" & "1111110000100111010101111101" & "00000001" & "10011100100010000010101001010011111110000100111010111000" & "10010100" & "1111111000010011101010111111" & "00000010" & "10011100100010000010101001010011111110000100111010110000" & "01001010" & "0111111100001001110101011111" & "00000000" & "10010011100100010000010101001010011111110000100111011000" & "10100101" & "0011111110000100111010110000" & "00000000" & "11001001110010001000001010100101001111111000010011101000" & "01010010" & "1001111111000010011101011000" & "00000000" & "11100100111001000100000101010010100111111100001001111000" & "10101001" & "0100111111100001001110101100" & "00000001" & "11100100111001000100000101010010100111111100001001101000" & "01010100" & "1010011111110000100111010110" & "00000000" & "10111001001110010001000001010100101001111111000010011000" & "00101010" & "0101001111111000010011101011" & "00000000" & "11011100100111001000100000101010010100111111100001011000" & "00010101" & "0010100111111100001001110101" & "00000001" & "11011100100111001000100000101010010100111111100001011000" & "00001010" & "1001010011111110000100111011" & "00000000" & "10110111001001110010001000001010100101001111111000011000" & "00000101" & "0100101001111111000010011101" & "00000000" & "11011011100100111001000100000101010010100111111100001000" & "10000010" & "1010010100111111100001001111" & "00000001" & "11011011100100111001000100000101010010100111111011111000" & "01000001" & "0101001010011111110000100111" & "00000010" & "11011011100100111001000100000101010010100111111100001000" & "00100000" & "1010100101001111111000010100" & "00000011" & "11011011100100111001000100000101010010100111111100100000" & "00010000" & "0101010010100111111100001010" & "00000100" & "11011011100100111001000100000101010010100111111010111000" & "10001000" & "0010101001010011111110000101"
 & "00000101" & "11011011100100111001000100000101010010100111111001101000" & "01000100" & "0001010100101001111111000010" & "00000000" & "10000011011011100100111001000100000101010010101000000000" & "00100010" & "0000101010010100111111100001" & "00000000" & "11000001101101110010011100100010000010101001010100001000" & "10010001" & "0000010101001010011111110001" & "00000001" & "11000001101101110010011100100010000010101001010011110000" & "11001000" & "1000001010100101001111111000" & "00000010" & "11000001101101110010011100100010000010101001010100001000" & "11100100" & "0100000101010010100111111100" & "00000000" & "10011000001101101110010011100100010000010101001010100000" & "01110010" & "0010000010101001010011111110" & "00000000" & "11001100000110110111001001110010001000001010100101010000" & "00111001" & "0001000001010100101001111111" & "00000000" & "11100110000011011011100100111001000100000101010010101000" & "10011100" & "1000100000101010010101000000" & "00000000" & "11110011000001101101110010011100100010000010101001001000" & "01001110" & "0100010000010101001010100000" & "00000000" & "11111001100000110110111001001110010001000001010100101000" & "00100111" & "0010001000001010100101010000" & "00000001" & "11111001100000110110111001001110010001000001010100101000" & "10010011" & "1001000100000101010010101000" & "00000000" & "10111110011000001101101110010011100100010000010101010000" & "11001001" & "1100100010000010101001010100" & "00000001" & "10111110011000001101101110010011100100010000010101011000" & "11100100" & "1110010001000001010100101010" & "00000010" & "10111110011000001101101110010011100100010000010101000000" & "01110010" & "0111001000100000101010010101" & "00000011" & "10111110011000001101101110010011100100010000010101110000" & "10111001" & "0011100100010000010101001010" & "00000000" & "10001011111001100000110110111001001110010001000001011000" & "11011100" & "1001110010001000001010100101" & "00000001" & "10001011111001100000110110111001001110010001000001010000" & "01101110" & "0100111001000100000101010011" & "00000000"
 & "10100010111110011000001101101110010011100100010000010000" & "10110111" & "0010011100100010000010101001" & "00000001" & "10100010111110011000001101101110010011100100010000011000" & "11011011" & "1001001110010001000001010101" & "00000010" & "10100010111110011000001101101110010011100100010000011000" & "01101101" & "1100100111001000100000101010" & "00000011" & "10100010111110011000001101101110010011100100010000011000" & "00110110" & "1110010011100100010000010101" & "00000100" & "10100010111110011000001101101110010011100100010000011000" & "00011011" & "0111001001110010001000001011" & "00000101" & "10100010111110011000001101101110010011100100010000011000" & "00001101" & "1011100100111001000100000101" & "00000110" & "10100010111110011000001101101110010011100100010000011000" & "00000110" & "1101110010011100100010000011" & "00000111" & "10100010111110011000001101101110010011100100010000011000" & "10000011" & "0110111001001110010001000001" & "00001000" & "10100010111110011000001101101110010011100101100001111000" & "11000001" & "1011011100100111001000100001" & "00001001" & "10100010111110011000001101101110010011100100010000011000" & "01100000" & "1101101110010011100100010000" & "00001010" & "10100010111110011000001101101110010011100100010000011000" & "00110000" & "0110110111001001110010001000" & "00001011" & "10100010111110011000001101101110010011100100010000011000" & "10011000" & "0011011011100100111001000100" & "00001100" & "10100010111110011000001101101110010011100100010000011000" & "11001100" & "0001101101110010011100100010" & "00001101" & "10100010111110011000001101101110010011100100010000011000" & "11100110" & "0000110110111001001110010001" & "00001110" & "10100010111110011000001101101110010011100100010000011000" & "11110011" & "0000011011011100100111001001" & "00001111" & "10100010111110011000001101101110010011100100010000011000" & "11111001" & "1000001101101110010011100100" & "00010000" & "10100010111110011000001101101110010011100100010000011000" & "01111100" & "1100000110110111001001110010" & "00010001" & "10100010111110011000001101101110001001011000010110111000"
 & "10111110" & "0110000011011011100100111001" & "00010010" & "10100010111110011000001101101110010011100100010000011000" & "01011111" & "0011000001101101110010011101" & "00010011" & "10100010111110011000001101101110011000101010001101001000" & "00101111" & "1001100000110110111001001110" & "00010100" & "10100010111110011000001101101110010011100100010000011000" & "00010111" & "1100110000011011011100100111" & "00010101" & "10100010111110011000001101101110010011100100010000011000" & "10001011" & "1110011000001101101110010100" & "00010110" & "10100010111110011000001101101110010011100100010000011000" & "01000101" & "1111001100000110110111001010" & "00010111" & "10100010111110011000001101101110010011100100010000011000" & "10100010" & "1111100110000011011011100101" & "00011000" & "10100010111110011000001101110000110110100010101000101000" & "01010001" & "0111110011000001101101110010" & "00011001" & "10100010111110011000001101101110010011100100010000011000" & "00101000" & "1011111001100000110110111001" & "00011010" & "10100010111110011000001101101110010011100100010000011000" & "00010100" & "0101111100110000011011011101" & "00011011" & "10100010111110011000001101101110010011100100010000011000" & "00001010" & "0010111110011000001101101110" & "00011100" & "10100010111110011000001101101110010011100100010000011000" & "00000101" & "0001011111001100000110110111" & "00011101" & "10100010111110011000001101101110010011100100010000011000" & "00000010" & "1000101111100110000011011100" & "00011110" & "10100010111110011000001101101110010011100100010000011000" & "00000001" & "0100010111110011000001101110" & "00011111" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "1010001011111001100000110111" & "00100000" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0101000101111100110000011011" & "00100001" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0010100010111110011000001110" & "00100010" & "10100010111110011000001101101110010011100100010000011000" & "00000000"
 & "0001010001011111001100000111" & "00100011" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000101000101111100110000011" & "00100100" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000010100010111110011000010" & "00100101" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000001010001011111001100001" & "00100110" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000101000101111100110000" & "00100111" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000010100010111110011000" & "00101000" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000001010001011111001100" & "00101001" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000000101000101111100110" & "00101010" & "10100010111110011000001101101110010011100100010000011000" & "00000000" & "0000000000010100010111110011" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
 & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
	loop36 : FOR i IN 0 TO 255 GENERATE
		loop37 : FOR j IN 0 TO 99 GENERATE
			wire_mux2_data_2d(i, j) <= wire_mux2_data(i*100+j);
		END GENERATE loop37;
	END GENERATE loop36;
	mux2 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 256,
		LPM_WIDTH => 100,
		LPM_WIDTHS => 8
	  )
	  PORT MAP ( 
		data => wire_mux2_data_2d,
		result => wire_mux2_result,
		sel => address
	  );

 END RTL; --coshw_altfp_sincos_srrt_koa


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altpriority_encoder_3e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END coshw_altpriority_encoder_3e8;

 ARCHITECTURE RTL OF coshw_altpriority_encoder_3e8 IS

 BEGIN

	q(0) <= ( data(1));
	zero <= (NOT (data(0) OR data(1)));

 END RTL; --coshw_altpriority_encoder_3e8


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=2 WIDTHAD=1 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altpriority_encoder_3v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0)
	 ); 
 END coshw_altpriority_encoder_3v7;

 ARCHITECTURE RTL OF coshw_altpriority_encoder_3v7 IS

 BEGIN

	q(0) <= ( data(1));

 END RTL; --coshw_altpriority_encoder_3v7

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altpriority_encoder_6v7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0)
	 ); 
 END coshw_altpriority_encoder_6v7;

 ARCHITECTURE RTL OF coshw_altpriority_encoder_6v7 IS

	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero12249w12250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero12251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_zero12249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_w_lg_w_lg_zero12251w12252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder10_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder9_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  coshw_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altpriority_encoder_3v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder10_w_lg_zero12249w & wire_altpriority_encoder10_w_lg_w_lg_zero12251w12252w);
	wire_altpriority_encoder10_w_lg_w_lg_zero12249w12250w(0) <= wire_altpriority_encoder10_w_lg_zero12249w(0) AND wire_altpriority_encoder10_q(0);
	wire_altpriority_encoder10_w_lg_zero12251w(0) <= wire_altpriority_encoder10_zero AND wire_altpriority_encoder9_q(0);
	wire_altpriority_encoder10_w_lg_zero12249w(0) <= NOT wire_altpriority_encoder10_zero;
	wire_altpriority_encoder10_w_lg_w_lg_zero12251w12252w(0) <= wire_altpriority_encoder10_w_lg_zero12251w(0) OR wire_altpriority_encoder10_w_lg_w_lg_zero12249w12250w(0);
	altpriority_encoder10 :  coshw_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder10_q,
		zero => wire_altpriority_encoder10_zero
	  );
	altpriority_encoder9 :  coshw_altpriority_encoder_3v7
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder9_q
	  );

 END RTL; --coshw_altpriority_encoder_6v7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=4 WIDTHAD=2 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altpriority_encoder_6e8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END coshw_altpriority_encoder_6e8;

 ARCHITECTURE RTL OF coshw_altpriority_encoder_6e8 IS

	 SIGNAL  wire_altpriority_encoder11_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder11_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero12267w12268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero12269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_zero12267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_w_lg_w_lg_zero12269w12270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_q	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder12_zero	:	STD_LOGIC;
	 COMPONENT  coshw_altpriority_encoder_3e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder12_w_lg_zero12267w & wire_altpriority_encoder12_w_lg_w_lg_zero12269w12270w);
	zero <= (wire_altpriority_encoder11_zero AND wire_altpriority_encoder12_zero);
	altpriority_encoder11 :  coshw_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(1 DOWNTO 0),
		q => wire_altpriority_encoder11_q,
		zero => wire_altpriority_encoder11_zero
	  );
	wire_altpriority_encoder12_w_lg_w_lg_zero12267w12268w(0) <= wire_altpriority_encoder12_w_lg_zero12267w(0) AND wire_altpriority_encoder12_q(0);
	wire_altpriority_encoder12_w_lg_zero12269w(0) <= wire_altpriority_encoder12_zero AND wire_altpriority_encoder11_q(0);
	wire_altpriority_encoder12_w_lg_zero12267w(0) <= NOT wire_altpriority_encoder12_zero;
	wire_altpriority_encoder12_w_lg_w_lg_zero12269w12270w(0) <= wire_altpriority_encoder12_w_lg_zero12269w(0) OR wire_altpriority_encoder12_w_lg_w_lg_zero12267w12268w(0);
	altpriority_encoder12 :  coshw_altpriority_encoder_3e8
	  PORT MAP ( 
		data => data(3 DOWNTO 2),
		q => wire_altpriority_encoder12_q,
		zero => wire_altpriority_encoder12_zero
	  );

 END RTL; --coshw_altpriority_encoder_6e8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altpriority_encoder_bv7 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END coshw_altpriority_encoder_bv7;

 ARCHITECTURE RTL OF coshw_altpriority_encoder_bv7 IS

	 SIGNAL  wire_altpriority_encoder7_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_w_lg_zero12240w12241w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_zero12242w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_zero12240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_w_lg_w_lg_zero12242w12243w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder8_zero	:	STD_LOGIC;
	 COMPONENT  coshw_altpriority_encoder_6v7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder8_w_lg_zero12240w & wire_altpriority_encoder8_w_lg_w_lg_zero12242w12243w);
	altpriority_encoder7 :  coshw_altpriority_encoder_6v7
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder7_q
	  );
	loop38 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder8_w_lg_w_lg_zero12240w12241w(i) <= wire_altpriority_encoder8_w_lg_zero12240w(0) AND wire_altpriority_encoder8_q(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder8_w_lg_zero12242w(i) <= wire_altpriority_encoder8_zero AND wire_altpriority_encoder7_q(i);
	END GENERATE loop39;
	wire_altpriority_encoder8_w_lg_zero12240w(0) <= NOT wire_altpriority_encoder8_zero;
	loop40 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder8_w_lg_w_lg_zero12242w12243w(i) <= wire_altpriority_encoder8_w_lg_zero12242w(i) OR wire_altpriority_encoder8_w_lg_w_lg_zero12240w12241w(i);
	END GENERATE loop40;
	altpriority_encoder8 :  coshw_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder8_q,
		zero => wire_altpriority_encoder8_zero
	  );

 END RTL; --coshw_altpriority_encoder_bv7


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=8 WIDTHAD=3 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altpriority_encoder_be8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END coshw_altpriority_encoder_be8;

 ARCHITECTURE RTL OF coshw_altpriority_encoder_be8 IS

	 SIGNAL  wire_altpriority_encoder13_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder13_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero12277w12278w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero12279w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_zero12277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_w_lg_w_lg_zero12279w12280w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_q	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder14_zero	:	STD_LOGIC;
	 COMPONENT  coshw_altpriority_encoder_6e8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder14_w_lg_zero12277w & wire_altpriority_encoder14_w_lg_w_lg_zero12279w12280w);
	zero <= (wire_altpriority_encoder13_zero AND wire_altpriority_encoder14_zero);
	altpriority_encoder13 :  coshw_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(3 DOWNTO 0),
		q => wire_altpriority_encoder13_q,
		zero => wire_altpriority_encoder13_zero
	  );
	loop41 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero12277w12278w(i) <= wire_altpriority_encoder14_w_lg_zero12277w(0) AND wire_altpriority_encoder14_q(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_zero12279w(i) <= wire_altpriority_encoder14_zero AND wire_altpriority_encoder13_q(i);
	END GENERATE loop42;
	wire_altpriority_encoder14_w_lg_zero12277w(0) <= NOT wire_altpriority_encoder14_zero;
	loop43 : FOR i IN 0 TO 1 GENERATE 
		wire_altpriority_encoder14_w_lg_w_lg_zero12279w12280w(i) <= wire_altpriority_encoder14_w_lg_zero12279w(i) OR wire_altpriority_encoder14_w_lg_w_lg_zero12277w12278w(i);
	END GENERATE loop43;
	altpriority_encoder14 :  coshw_altpriority_encoder_6e8
	  PORT MAP ( 
		data => data(7 DOWNTO 4),
		q => wire_altpriority_encoder14_q,
		zero => wire_altpriority_encoder14_zero
	  );

 END RTL; --coshw_altpriority_encoder_be8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altpriority_encoder_r08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0)
	 ); 
 END coshw_altpriority_encoder_r08;

 ARCHITECTURE RTL OF coshw_altpriority_encoder_r08 IS

	 SIGNAL  wire_altpriority_encoder5_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_w_lg_w_lg_zero12231w12232w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_w_lg_zero12233w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_w_lg_zero12231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_w_lg_w_lg_zero12233w12234w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder6_zero	:	STD_LOGIC;
	 COMPONENT  coshw_altpriority_encoder_bv7
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder6_w_lg_zero12231w & wire_altpriority_encoder6_w_lg_w_lg_zero12233w12234w);
	altpriority_encoder5 :  coshw_altpriority_encoder_bv7
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder5_q
	  );
	loop44 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder6_w_lg_w_lg_zero12231w12232w(i) <= wire_altpriority_encoder6_w_lg_zero12231w(0) AND wire_altpriority_encoder6_q(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder6_w_lg_zero12233w(i) <= wire_altpriority_encoder6_zero AND wire_altpriority_encoder5_q(i);
	END GENERATE loop45;
	wire_altpriority_encoder6_w_lg_zero12231w(0) <= NOT wire_altpriority_encoder6_zero;
	loop46 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder6_w_lg_w_lg_zero12233w12234w(i) <= wire_altpriority_encoder6_w_lg_zero12233w(i) OR wire_altpriority_encoder6_w_lg_w_lg_zero12231w12232w(i);
	END GENERATE loop46;
	altpriority_encoder6 :  coshw_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder6_q,
		zero => wire_altpriority_encoder6_zero
	  );

 END RTL; --coshw_altpriority_encoder_r08


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=16 WIDTHAD=4 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altpriority_encoder_rf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END coshw_altpriority_encoder_rf8;

 ARCHITECTURE RTL OF coshw_altpriority_encoder_rf8 IS

	 SIGNAL  wire_altpriority_encoder15_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder15_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero12287w12288w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero12289w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_zero12287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_w_lg_w_lg_zero12289w12290w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder16_zero	:	STD_LOGIC;
	 COMPONENT  coshw_altpriority_encoder_be8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder16_w_lg_zero12287w & wire_altpriority_encoder16_w_lg_w_lg_zero12289w12290w);
	zero <= (wire_altpriority_encoder15_zero AND wire_altpriority_encoder16_zero);
	altpriority_encoder15 :  coshw_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(7 DOWNTO 0),
		q => wire_altpriority_encoder15_q,
		zero => wire_altpriority_encoder15_zero
	  );
	loop47 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder16_w_lg_w_lg_zero12287w12288w(i) <= wire_altpriority_encoder16_w_lg_zero12287w(0) AND wire_altpriority_encoder16_q(i);
	END GENERATE loop47;
	loop48 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder16_w_lg_zero12289w(i) <= wire_altpriority_encoder16_zero AND wire_altpriority_encoder15_q(i);
	END GENERATE loop48;
	wire_altpriority_encoder16_w_lg_zero12287w(0) <= NOT wire_altpriority_encoder16_zero;
	loop49 : FOR i IN 0 TO 2 GENERATE 
		wire_altpriority_encoder16_w_lg_w_lg_zero12289w12290w(i) <= wire_altpriority_encoder16_w_lg_zero12289w(i) OR wire_altpriority_encoder16_w_lg_w_lg_zero12287w12288w(i);
	END GENERATE loop49;
	altpriority_encoder16 :  coshw_altpriority_encoder_be8
	  PORT MAP ( 
		data => data(15 DOWNTO 8),
		q => wire_altpriority_encoder16_q,
		zero => wire_altpriority_encoder16_zero
	  );

 END RTL; --coshw_altpriority_encoder_rf8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altpriority_encoder_qb6 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END coshw_altpriority_encoder_qb6;

 ARCHITECTURE RTL OF coshw_altpriority_encoder_qb6 IS

	 SIGNAL  wire_altpriority_encoder3_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_w_lg_w_lg_zero12222w12223w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_w_lg_zero12224w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_w_lg_zero12222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_w_lg_w_lg_zero12224w12225w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder4_zero	:	STD_LOGIC;
	 COMPONENT  coshw_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder4_w_lg_zero12222w & wire_altpriority_encoder4_w_lg_w_lg_zero12224w12225w);
	altpriority_encoder3 :  coshw_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder3_q
	  );
	loop50 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder4_w_lg_w_lg_zero12222w12223w(i) <= wire_altpriority_encoder4_w_lg_zero12222w(0) AND wire_altpriority_encoder4_q(i);
	END GENERATE loop50;
	loop51 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder4_w_lg_zero12224w(i) <= wire_altpriority_encoder4_zero AND wire_altpriority_encoder3_q(i);
	END GENERATE loop51;
	wire_altpriority_encoder4_w_lg_zero12222w(0) <= NOT wire_altpriority_encoder4_zero;
	loop52 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder4_w_lg_w_lg_zero12224w12225w(i) <= wire_altpriority_encoder4_w_lg_zero12224w(i) OR wire_altpriority_encoder4_w_lg_w_lg_zero12222w12223w(i);
	END GENERATE loop52;
	altpriority_encoder4 :  coshw_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder4_q,
		zero => wire_altpriority_encoder4_zero
	  );

 END RTL; --coshw_altpriority_encoder_qb6

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 8 lpm_clshift 2 lpm_mult 1 lpm_mux 1 reg 780 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_range_b6c IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 circle	:	OUT  STD_LOGIC_VECTOR (35 DOWNTO 0);
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0) := (OTHERS => '0');
		 negcircle	:	OUT  STD_LOGIC_VECTOR (35 DOWNTO 0)
	 ); 
 END coshw_altfp_sincos_range_b6c;

 ARCHITECTURE RTL OF coshw_altfp_sincos_range_b6c IS

	 SIGNAL  wire_fp_range_table1_basefraction	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_fp_range_table1_incexponent	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_fp_range_table1_incmantissa	:	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  wire_clz23_data	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_clz23_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL	 basefractiondelff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 basefractionff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_0	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_1	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_2	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_3	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_4	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 cbfd_5	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 circleff	:	STD_LOGIC_VECTOR(36 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponentff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 incexponentff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 incmantissaff	:	STD_LOGIC_VECTOR(55 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 leadff	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissadelff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissaff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissamultiplierff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 multipliernormff	:	STD_LOGIC_VECTOR(77 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 negbasefractiondelff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 negcircleff	:	STD_LOGIC_VECTOR(36 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 negrangeexponentff4	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 negrangeexponentff5	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_negrangeexponentff5_w_lg_w_lg_w_q_range10692w10696w10697w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_lg_w_q_range10692w10694w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_lg_w_q_range10692w10696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_q_range10693w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_q_range10692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rangeexponentff_0	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_1	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_2	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_3	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_4	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rangeexponentff_5	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rangeexponentff_5_w_q_range10695w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL	 rotateff	:	STD_LOGIC_VECTOR(77 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rotateff_w_lg_w_q_range10709w10710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10713w10714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10716w10717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10719w10720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10722w10723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10725w10726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10728w10729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10731w10732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10734w10735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10737w10738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10740w10741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10743w10744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10746w10747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10749w10750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10752w10753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10755w10756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10758w10759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10761w10762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10764w10765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10767w10768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10770w10771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10773w10774w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10776w10777w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10779w10780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10782w10783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10785w10786w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10788w10789w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10791w10792w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10794w10795w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10797w10798w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10800w10801w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10803w10804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10806w10807w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10809w10810w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10812w10813w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_lg_w_q_range10815w10816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10782w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10785w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10791w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10794w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10797w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10803w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10806w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10809w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10812w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rotateff_w_q_range10815w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 tableaddressff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_circle_add_dataa	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_circle_add_datab	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_circle_add_result	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_exponent_adjust_sub_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_exponent_adjust_sub_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_negbasedractiondel_sub_dataa	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_negbasedractiondel_sub_result	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_negcircle_add_dataa	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_negcircle_add_datab	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_negcircle_add_result	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_negrangeexponent_sub4_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_negrangeexponent_sub4_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_negrangeexponent_sub5_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_negrangeexponent_sub5_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rangeexponent_sub1_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rangeexponent_sub1_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rangeexponent_sub5_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rangeexponent_sub5_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_csftin_result	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_fp_lsft_rsft78_distance	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_negrangeexponentff5_w_lg_w_lg_w_lg_w_q_range10692w10696w10697w10698w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_fp_lsft_rsft78_result	:	STD_LOGIC_VECTOR (77 DOWNTO 0);
	 SIGNAL  wire_mult23x56_result	:	STD_LOGIC_VECTOR (78 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10301w10302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10349w10353w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10349w10350w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10354w10358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10354w10355w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10359w10363w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10359w10360w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10364w10368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10364w10365w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10369w10373w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10369w10370w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10374w10378w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10374w10375w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10379w10383w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10379w10380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10384w10388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10384w10385w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10389w10393w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10389w10390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10394w10398w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10394w10395w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10303w10308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10303w10304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10399w10403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10399w10400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10404w10408w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10404w10405w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10409w10413w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10409w10410w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10414w10418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10414w10415w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10419w10423w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10419w10420w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10424w10428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10424w10425w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10429w10433w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10429w10430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10434w10438w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10434w10435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10439w10443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10439w10440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10444w10448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10444w10445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10309w10313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10309w10310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10449w10453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10449w10450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10454w10458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10454w10455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10459w10463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10459w10460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10464w10468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10464w10465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10469w10473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10469w10470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10474w10478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10474w10475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10479w10483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10479w10480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10484w10488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10484w10485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10489w10493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10489w10490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10494w10498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10494w10495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10314w10318w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10314w10315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10499w10503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10499w10500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10504w10508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10504w10505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10509w10513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10509w10510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10514w10518w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10514w10515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10519w10523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10519w10520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10524w10528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10524w10525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10529w10533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10529w10530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10534w10538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10534w10535w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10539w10543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10539w10540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10544w10548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10544w10545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10319w10323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10319w10320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10549w10553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10549w10550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10554w10558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10554w10555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10559w10563w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10559w10560w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10564w10568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10564w10565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10569w10573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10569w10570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10574w10578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10574w10575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10579w10583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10579w10580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10584w10588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10584w10585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10589w10593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10589w10590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10594w10598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10594w10595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10324w10328w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10324w10325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10599w10603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10599w10600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10604w10608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10604w10605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10609w10613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10609w10610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10614w10618w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10614w10615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10619w10623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10619w10620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10624w10628w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10624w10625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10629w10633w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10629w10630w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10634w10638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10634w10635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10639w10643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10639w10640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10644w10648w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10644w10645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10329w10333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10329w10330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10649w10653w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10649w10650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10654w10658w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10654w10655w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10659w10663w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10659w10660w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10664w10668w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10664w10665w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10669w10673w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10669w10670w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10674w10678w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10674w10675w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10679w10683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10679w10680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10684w10688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10684w10685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10334w10338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10334w10335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10339w10343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10339w10340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10344w10348w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10344w10345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10371w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10376w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10381w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10386w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10396w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10406w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10416w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10421w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10426w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10431w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10316w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10561w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10326w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10621w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10626w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10631w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10636w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10646w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10656w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10661w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10666w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10671w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10336w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w10346w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  basefractiondelnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  basefractionnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  circlenode_w :	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  const_23_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  incexponentnode_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  incmantissanode_w :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  leadnode_w :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  mantissaexponentnode_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  mantissamultipliernode_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  multipliernode_w :	STD_LOGIC_VECTOR (78 DOWNTO 0);
	 SIGNAL  multipliernormnode_w :	STD_LOGIC_VECTOR (77 DOWNTO 0);
	 SIGNAL  negbasefractiondelnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  negcirclenode_w :	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  negrotatenode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  rotatenode_w :	STD_LOGIC_VECTOR (77 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_data_range10271w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_data_range10272w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10354w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10369w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10374w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10379w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10384w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10389w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10399w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10409w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10419w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10424w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10429w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10434w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10319w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10559w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10634w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10639w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10654w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10659w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10664w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10669w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10679w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_w_multipliernode_w_range10344w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  coshw_altfp_sincos_srrt_koa
	 PORT
	 ( 
		address	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		basefraction	:	OUT  STD_LOGIC_VECTOR(35 DOWNTO 0);
		incexponent	:	OUT  STD_LOGIC_VECTOR(7 DOWNTO 0);
		incmantissa	:	OUT  STD_LOGIC_VECTOR(55 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altpriority_encoder_qb6
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_clshift
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_SHIFTTYPE	:	STRING := "LOGICAL";
		LPM_WIDTH	:	NATURAL;
		LPM_WIDTHDIST	:	NATURAL;
		lpm_type	:	STRING := "lpm_clshift"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		direction	:	IN STD_LOGIC := '0';
		distance	:	IN STD_LOGIC_VECTOR(LPM_WIDTHDIST-1 DOWNTO 0);
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		underflow	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_vcc <= '1';
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10301w10302w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10301w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10349w10353w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10349w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10349w10350w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10349w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10354w10358w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10354w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10354w10355w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10354w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10359w10363w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10359w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10359w10360w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10359w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10364w10368w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10364w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10364w10365w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10364w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10369w10373w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10369w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10369w10370w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10369w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10374w10378w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10374w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10374w10375w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10374w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10379w10383w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10379w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10379w10380w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10379w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10384w10388w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10384w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10384w10385w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10384w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10389w10393w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10389w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10389w10390w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10389w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10394w10398w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10394w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10394w10395w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10394w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10303w10308w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10303w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10303w10304w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10303w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10399w10403w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10399w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10399w10400w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10399w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10404w10408w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10404w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10404w10405w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10404w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10409w10413w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10409w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10409w10410w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10409w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10414w10418w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10414w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10414w10415w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10414w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10419w10423w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10419w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10419w10420w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10419w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10424w10428w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10424w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10424w10425w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10424w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10429w10433w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10429w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10429w10430w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10429w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10434w10438w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10434w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10434w10435w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10434w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10439w10443w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10439w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10439w10440w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10439w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10444w10448w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10444w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10444w10445w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10444w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10309w10313w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10309w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10309w10310w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10309w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10449w10453w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10449w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10449w10450w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10449w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10454w10458w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10454w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10454w10455w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10454w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10459w10463w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10459w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10459w10460w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10459w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10464w10468w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10464w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10464w10465w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10464w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10469w10473w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10469w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10469w10470w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10469w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10474w10478w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10474w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10474w10475w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10474w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10479w10483w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10479w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10479w10480w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10479w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10484w10488w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10484w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10484w10485w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10484w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10489w10493w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10489w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10489w10490w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10489w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10494w10498w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10494w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10494w10495w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10494w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10314w10318w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10314w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10314w10315w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10314w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10499w10503w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10499w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10499w10500w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10499w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10504w10508w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10504w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10504w10505w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10504w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10509w10513w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10509w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10509w10510w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10509w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10514w10518w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10514w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10514w10515w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10514w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10519w10523w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10519w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10519w10520w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10519w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10524w10528w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10524w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10524w10525w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10524w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10529w10533w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10529w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10529w10530w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10529w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10534w10538w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10534w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10534w10535w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10534w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10539w10543w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10539w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10539w10540w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10539w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10544w10548w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10544w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10544w10545w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10544w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10319w10323w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10319w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10319w10320w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10319w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10549w10553w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10549w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10549w10550w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10549w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10554w10558w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10554w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10554w10555w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10554w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10559w10563w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10559w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10559w10560w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10559w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10564w10568w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10564w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10564w10565w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10564w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10569w10573w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10569w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10569w10570w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10569w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10574w10578w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10574w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10574w10575w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10574w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10579w10583w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10579w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10579w10580w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10579w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10584w10588w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10584w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10584w10585w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10584w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10589w10593w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10589w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10589w10590w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10589w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10594w10598w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10594w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10594w10595w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10594w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10324w10328w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10324w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10324w10325w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10324w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10599w10603w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10599w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10599w10600w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10599w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10604w10608w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10604w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10604w10605w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10604w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10609w10613w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10609w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10609w10610w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10609w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10614w10618w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10614w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10614w10615w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10614w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10619w10623w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10619w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10619w10620w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10619w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10624w10628w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10624w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10624w10625w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10624w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10629w10633w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10629w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10629w10630w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10629w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10634w10638w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10634w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10634w10635w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10634w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10639w10643w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10639w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10639w10640w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10639w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10644w10648w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10644w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10644w10645w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10644w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10329w10333w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10329w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10329w10330w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10329w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10649w10653w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10649w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10649w10650w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10649w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10654w10658w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10654w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10654w10655w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10654w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10659w10663w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10659w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10659w10660w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10659w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10664w10668w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10664w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10664w10665w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10664w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10669w10673w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10669w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10669w10670w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10669w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10674w10678w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10674w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10674w10675w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10674w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10679w10683w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10679w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10679w10680w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10679w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10684w10688w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10684w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10684w10685w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10684w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10689w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10280w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10334w10338w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10334w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10334w10335w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10334w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10339w10343w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10339w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10339w10340w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10339w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10344w10348w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10344w(0) AND wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10344w10345w(0) <= wire_crr_fp_range1_w_multipliernode_w_range10344w(0) AND wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w(0) <= NOT wire_crr_fp_range1_w_multipliernode_w_range10280w(0);
	wire_crr_fp_range1_w10351w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10349w10350w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10344w10348w(0);
	wire_crr_fp_range1_w10356w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10354w10355w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10349w10353w(0);
	wire_crr_fp_range1_w10361w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10359w10360w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10354w10358w(0);
	wire_crr_fp_range1_w10366w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10364w10365w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10359w10363w(0);
	wire_crr_fp_range1_w10371w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10369w10370w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10364w10368w(0);
	wire_crr_fp_range1_w10376w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10374w10375w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10369w10373w(0);
	wire_crr_fp_range1_w10381w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10379w10380w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10374w10378w(0);
	wire_crr_fp_range1_w10386w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10384w10385w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10379w10383w(0);
	wire_crr_fp_range1_w10391w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10389w10390w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10384w10388w(0);
	wire_crr_fp_range1_w10396w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10394w10395w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10389w10393w(0);
	wire_crr_fp_range1_w10305w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10303w10304w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10301w10302w(0);
	wire_crr_fp_range1_w10401w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10399w10400w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10394w10398w(0);
	wire_crr_fp_range1_w10406w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10404w10405w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10399w10403w(0);
	wire_crr_fp_range1_w10411w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10409w10410w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10404w10408w(0);
	wire_crr_fp_range1_w10416w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10414w10415w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10409w10413w(0);
	wire_crr_fp_range1_w10421w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10419w10420w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10414w10418w(0);
	wire_crr_fp_range1_w10426w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10424w10425w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10419w10423w(0);
	wire_crr_fp_range1_w10431w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10429w10430w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10424w10428w(0);
	wire_crr_fp_range1_w10436w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10434w10435w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10429w10433w(0);
	wire_crr_fp_range1_w10441w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10439w10440w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10434w10438w(0);
	wire_crr_fp_range1_w10446w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10444w10445w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10439w10443w(0);
	wire_crr_fp_range1_w10311w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10309w10310w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10303w10308w(0);
	wire_crr_fp_range1_w10451w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10449w10450w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10444w10448w(0);
	wire_crr_fp_range1_w10456w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10454w10455w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10449w10453w(0);
	wire_crr_fp_range1_w10461w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10459w10460w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10454w10458w(0);
	wire_crr_fp_range1_w10466w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10464w10465w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10459w10463w(0);
	wire_crr_fp_range1_w10471w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10469w10470w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10464w10468w(0);
	wire_crr_fp_range1_w10476w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10474w10475w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10469w10473w(0);
	wire_crr_fp_range1_w10481w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10479w10480w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10474w10478w(0);
	wire_crr_fp_range1_w10486w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10484w10485w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10479w10483w(0);
	wire_crr_fp_range1_w10491w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10489w10490w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10484w10488w(0);
	wire_crr_fp_range1_w10496w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10494w10495w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10489w10493w(0);
	wire_crr_fp_range1_w10316w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10314w10315w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10309w10313w(0);
	wire_crr_fp_range1_w10501w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10499w10500w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10494w10498w(0);
	wire_crr_fp_range1_w10506w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10504w10505w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10499w10503w(0);
	wire_crr_fp_range1_w10511w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10509w10510w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10504w10508w(0);
	wire_crr_fp_range1_w10516w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10514w10515w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10509w10513w(0);
	wire_crr_fp_range1_w10521w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10519w10520w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10514w10518w(0);
	wire_crr_fp_range1_w10526w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10524w10525w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10519w10523w(0);
	wire_crr_fp_range1_w10531w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10529w10530w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10524w10528w(0);
	wire_crr_fp_range1_w10536w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10534w10535w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10529w10533w(0);
	wire_crr_fp_range1_w10541w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10539w10540w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10534w10538w(0);
	wire_crr_fp_range1_w10546w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10544w10545w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10539w10543w(0);
	wire_crr_fp_range1_w10321w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10319w10320w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10314w10318w(0);
	wire_crr_fp_range1_w10551w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10549w10550w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10544w10548w(0);
	wire_crr_fp_range1_w10556w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10554w10555w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10549w10553w(0);
	wire_crr_fp_range1_w10561w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10559w10560w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10554w10558w(0);
	wire_crr_fp_range1_w10566w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10564w10565w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10559w10563w(0);
	wire_crr_fp_range1_w10571w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10569w10570w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10564w10568w(0);
	wire_crr_fp_range1_w10576w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10574w10575w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10569w10573w(0);
	wire_crr_fp_range1_w10581w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10579w10580w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10574w10578w(0);
	wire_crr_fp_range1_w10586w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10584w10585w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10579w10583w(0);
	wire_crr_fp_range1_w10591w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10589w10590w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10584w10588w(0);
	wire_crr_fp_range1_w10596w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10594w10595w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10589w10593w(0);
	wire_crr_fp_range1_w10326w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10324w10325w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10319w10323w(0);
	wire_crr_fp_range1_w10601w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10599w10600w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10594w10598w(0);
	wire_crr_fp_range1_w10606w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10604w10605w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10599w10603w(0);
	wire_crr_fp_range1_w10611w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10609w10610w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10604w10608w(0);
	wire_crr_fp_range1_w10616w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10614w10615w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10609w10613w(0);
	wire_crr_fp_range1_w10621w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10619w10620w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10614w10618w(0);
	wire_crr_fp_range1_w10626w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10624w10625w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10619w10623w(0);
	wire_crr_fp_range1_w10631w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10629w10630w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10624w10628w(0);
	wire_crr_fp_range1_w10636w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10634w10635w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10629w10633w(0);
	wire_crr_fp_range1_w10641w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10639w10640w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10634w10638w(0);
	wire_crr_fp_range1_w10646w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10644w10645w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10639w10643w(0);
	wire_crr_fp_range1_w10331w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10329w10330w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10324w10328w(0);
	wire_crr_fp_range1_w10651w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10649w10650w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10644w10648w(0);
	wire_crr_fp_range1_w10656w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10654w10655w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10649w10653w(0);
	wire_crr_fp_range1_w10661w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10659w10660w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10654w10658w(0);
	wire_crr_fp_range1_w10666w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10664w10665w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10659w10663w(0);
	wire_crr_fp_range1_w10671w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10669w10670w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10664w10668w(0);
	wire_crr_fp_range1_w10676w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10674w10675w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10669w10673w(0);
	wire_crr_fp_range1_w10681w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10679w10680w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10674w10678w(0);
	wire_crr_fp_range1_w10686w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10684w10685w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10679w10683w(0);
	wire_crr_fp_range1_w10690w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10689w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10684w10688w(0);
	wire_crr_fp_range1_w10336w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10334w10335w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10329w10333w(0);
	wire_crr_fp_range1_w10341w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10339w10340w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10334w10338w(0);
	wire_crr_fp_range1_w10346w(0) <= wire_crr_fp_range1_w_lg_w_multipliernode_w_range10344w10345w(0) OR wire_crr_fp_range1_w_lg_w_multipliernode_w_range10339w10343w(0);
	basefractiondelnode_w <= cbfd_5;
	basefractionnode_w <= wire_fp_range_table1_basefraction;
	circle <= circleff(35 DOWNTO 0);
	circlenode_w <= wire_circle_add_result;
	const_23_w <= "000010111";
	incexponentnode_w <= wire_fp_range_table1_incexponent;
	incmantissanode_w <= wire_fp_range_table1_incmantissa;
	leadnode_w <= (NOT wire_clz23_q);
	mantissaexponentnode_w <= wire_exponent_adjust_sub_result;
	mantissamultipliernode_w <= wire_csftin_result;
	multipliernode_w <= wire_mult23x56_result;
	multipliernormnode_w <= ( wire_crr_fp_range1_w10690w & wire_crr_fp_range1_w10686w & wire_crr_fp_range1_w10681w & wire_crr_fp_range1_w10676w & wire_crr_fp_range1_w10671w & wire_crr_fp_range1_w10666w & wire_crr_fp_range1_w10661w & wire_crr_fp_range1_w10656w & wire_crr_fp_range1_w10651w & wire_crr_fp_range1_w10646w & wire_crr_fp_range1_w10641w & wire_crr_fp_range1_w10636w & wire_crr_fp_range1_w10631w & wire_crr_fp_range1_w10626w & wire_crr_fp_range1_w10621w & wire_crr_fp_range1_w10616w & wire_crr_fp_range1_w10611w & wire_crr_fp_range1_w10606w & wire_crr_fp_range1_w10601w & wire_crr_fp_range1_w10596w & wire_crr_fp_range1_w10591w & wire_crr_fp_range1_w10586w & wire_crr_fp_range1_w10581w & wire_crr_fp_range1_w10576w & wire_crr_fp_range1_w10571w & wire_crr_fp_range1_w10566w & wire_crr_fp_range1_w10561w & wire_crr_fp_range1_w10556w & wire_crr_fp_range1_w10551w & wire_crr_fp_range1_w10546w & wire_crr_fp_range1_w10541w & wire_crr_fp_range1_w10536w & wire_crr_fp_range1_w10531w & wire_crr_fp_range1_w10526w & wire_crr_fp_range1_w10521w & wire_crr_fp_range1_w10516w & wire_crr_fp_range1_w10511w & wire_crr_fp_range1_w10506w & wire_crr_fp_range1_w10501w & wire_crr_fp_range1_w10496w & wire_crr_fp_range1_w10491w & wire_crr_fp_range1_w10486w & wire_crr_fp_range1_w10481w & wire_crr_fp_range1_w10476w & wire_crr_fp_range1_w10471w & wire_crr_fp_range1_w10466w & wire_crr_fp_range1_w10461w & wire_crr_fp_range1_w10456w & wire_crr_fp_range1_w10451w & wire_crr_fp_range1_w10446w & wire_crr_fp_range1_w10441w & wire_crr_fp_range1_w10436w & wire_crr_fp_range1_w10431w & wire_crr_fp_range1_w10426w & wire_crr_fp_range1_w10421w & wire_crr_fp_range1_w10416w & wire_crr_fp_range1_w10411w & wire_crr_fp_range1_w10406w & wire_crr_fp_range1_w10401w & wire_crr_fp_range1_w10396w & wire_crr_fp_range1_w10391w & wire_crr_fp_range1_w10386w & wire_crr_fp_range1_w10381w & wire_crr_fp_range1_w10376w & wire_crr_fp_range1_w10371w & wire_crr_fp_range1_w10366w & wire_crr_fp_range1_w10361w & wire_crr_fp_range1_w10356w & wire_crr_fp_range1_w10351w & wire_crr_fp_range1_w10346w
 & wire_crr_fp_range1_w10341w & wire_crr_fp_range1_w10336w & wire_crr_fp_range1_w10331w & wire_crr_fp_range1_w10326w & wire_crr_fp_range1_w10321w & wire_crr_fp_range1_w10316w & wire_crr_fp_range1_w10311w & wire_crr_fp_range1_w10305w);
	negbasefractiondelnode_w <= wire_negbasedractiondel_sub_result;
	negcircle <= negcircleff(35 DOWNTO 0);
	negcirclenode_w <= wire_negcircle_add_result;
	negrotatenode_w <= ( wire_rotateff_w_lg_w_q_range10815w10816w & wire_rotateff_w_lg_w_q_range10812w10813w & wire_rotateff_w_lg_w_q_range10809w10810w & wire_rotateff_w_lg_w_q_range10806w10807w & wire_rotateff_w_lg_w_q_range10803w10804w & wire_rotateff_w_lg_w_q_range10800w10801w & wire_rotateff_w_lg_w_q_range10797w10798w & wire_rotateff_w_lg_w_q_range10794w10795w & wire_rotateff_w_lg_w_q_range10791w10792w & wire_rotateff_w_lg_w_q_range10788w10789w & wire_rotateff_w_lg_w_q_range10785w10786w & wire_rotateff_w_lg_w_q_range10782w10783w & wire_rotateff_w_lg_w_q_range10779w10780w & wire_rotateff_w_lg_w_q_range10776w10777w & wire_rotateff_w_lg_w_q_range10773w10774w & wire_rotateff_w_lg_w_q_range10770w10771w & wire_rotateff_w_lg_w_q_range10767w10768w & wire_rotateff_w_lg_w_q_range10764w10765w & wire_rotateff_w_lg_w_q_range10761w10762w & wire_rotateff_w_lg_w_q_range10758w10759w & wire_rotateff_w_lg_w_q_range10755w10756w & wire_rotateff_w_lg_w_q_range10752w10753w & wire_rotateff_w_lg_w_q_range10749w10750w & wire_rotateff_w_lg_w_q_range10746w10747w & wire_rotateff_w_lg_w_q_range10743w10744w & wire_rotateff_w_lg_w_q_range10740w10741w & wire_rotateff_w_lg_w_q_range10737w10738w & wire_rotateff_w_lg_w_q_range10734w10735w & wire_rotateff_w_lg_w_q_range10731w10732w & wire_rotateff_w_lg_w_q_range10728w10729w & wire_rotateff_w_lg_w_q_range10725w10726w & wire_rotateff_w_lg_w_q_range10722w10723w & wire_rotateff_w_lg_w_q_range10719w10720w & wire_rotateff_w_lg_w_q_range10716w10717w & wire_rotateff_w_lg_w_q_range10713w10714w & wire_rotateff_w_lg_w_q_range10709w10710w);
	rotatenode_w <= wire_fp_lsft_rsft78_result;
	wire_crr_fp_range1_w_data_range10271w <= data(22 DOWNTO 0);
	wire_crr_fp_range1_w_data_range10272w <= data(30 DOWNTO 23);
	wire_crr_fp_range1_w_multipliernode_w_range10301w(0) <= multipliernode_w(0);
	wire_crr_fp_range1_w_multipliernode_w_range10349w(0) <= multipliernode_w(10);
	wire_crr_fp_range1_w_multipliernode_w_range10354w(0) <= multipliernode_w(11);
	wire_crr_fp_range1_w_multipliernode_w_range10359w(0) <= multipliernode_w(12);
	wire_crr_fp_range1_w_multipliernode_w_range10364w(0) <= multipliernode_w(13);
	wire_crr_fp_range1_w_multipliernode_w_range10369w(0) <= multipliernode_w(14);
	wire_crr_fp_range1_w_multipliernode_w_range10374w(0) <= multipliernode_w(15);
	wire_crr_fp_range1_w_multipliernode_w_range10379w(0) <= multipliernode_w(16);
	wire_crr_fp_range1_w_multipliernode_w_range10384w(0) <= multipliernode_w(17);
	wire_crr_fp_range1_w_multipliernode_w_range10389w(0) <= multipliernode_w(18);
	wire_crr_fp_range1_w_multipliernode_w_range10394w(0) <= multipliernode_w(19);
	wire_crr_fp_range1_w_multipliernode_w_range10303w(0) <= multipliernode_w(1);
	wire_crr_fp_range1_w_multipliernode_w_range10399w(0) <= multipliernode_w(20);
	wire_crr_fp_range1_w_multipliernode_w_range10404w(0) <= multipliernode_w(21);
	wire_crr_fp_range1_w_multipliernode_w_range10409w(0) <= multipliernode_w(22);
	wire_crr_fp_range1_w_multipliernode_w_range10414w(0) <= multipliernode_w(23);
	wire_crr_fp_range1_w_multipliernode_w_range10419w(0) <= multipliernode_w(24);
	wire_crr_fp_range1_w_multipliernode_w_range10424w(0) <= multipliernode_w(25);
	wire_crr_fp_range1_w_multipliernode_w_range10429w(0) <= multipliernode_w(26);
	wire_crr_fp_range1_w_multipliernode_w_range10434w(0) <= multipliernode_w(27);
	wire_crr_fp_range1_w_multipliernode_w_range10439w(0) <= multipliernode_w(28);
	wire_crr_fp_range1_w_multipliernode_w_range10444w(0) <= multipliernode_w(29);
	wire_crr_fp_range1_w_multipliernode_w_range10309w(0) <= multipliernode_w(2);
	wire_crr_fp_range1_w_multipliernode_w_range10449w(0) <= multipliernode_w(30);
	wire_crr_fp_range1_w_multipliernode_w_range10454w(0) <= multipliernode_w(31);
	wire_crr_fp_range1_w_multipliernode_w_range10459w(0) <= multipliernode_w(32);
	wire_crr_fp_range1_w_multipliernode_w_range10464w(0) <= multipliernode_w(33);
	wire_crr_fp_range1_w_multipliernode_w_range10469w(0) <= multipliernode_w(34);
	wire_crr_fp_range1_w_multipliernode_w_range10474w(0) <= multipliernode_w(35);
	wire_crr_fp_range1_w_multipliernode_w_range10479w(0) <= multipliernode_w(36);
	wire_crr_fp_range1_w_multipliernode_w_range10484w(0) <= multipliernode_w(37);
	wire_crr_fp_range1_w_multipliernode_w_range10489w(0) <= multipliernode_w(38);
	wire_crr_fp_range1_w_multipliernode_w_range10494w(0) <= multipliernode_w(39);
	wire_crr_fp_range1_w_multipliernode_w_range10314w(0) <= multipliernode_w(3);
	wire_crr_fp_range1_w_multipliernode_w_range10499w(0) <= multipliernode_w(40);
	wire_crr_fp_range1_w_multipliernode_w_range10504w(0) <= multipliernode_w(41);
	wire_crr_fp_range1_w_multipliernode_w_range10509w(0) <= multipliernode_w(42);
	wire_crr_fp_range1_w_multipliernode_w_range10514w(0) <= multipliernode_w(43);
	wire_crr_fp_range1_w_multipliernode_w_range10519w(0) <= multipliernode_w(44);
	wire_crr_fp_range1_w_multipliernode_w_range10524w(0) <= multipliernode_w(45);
	wire_crr_fp_range1_w_multipliernode_w_range10529w(0) <= multipliernode_w(46);
	wire_crr_fp_range1_w_multipliernode_w_range10534w(0) <= multipliernode_w(47);
	wire_crr_fp_range1_w_multipliernode_w_range10539w(0) <= multipliernode_w(48);
	wire_crr_fp_range1_w_multipliernode_w_range10544w(0) <= multipliernode_w(49);
	wire_crr_fp_range1_w_multipliernode_w_range10319w(0) <= multipliernode_w(4);
	wire_crr_fp_range1_w_multipliernode_w_range10549w(0) <= multipliernode_w(50);
	wire_crr_fp_range1_w_multipliernode_w_range10554w(0) <= multipliernode_w(51);
	wire_crr_fp_range1_w_multipliernode_w_range10559w(0) <= multipliernode_w(52);
	wire_crr_fp_range1_w_multipliernode_w_range10564w(0) <= multipliernode_w(53);
	wire_crr_fp_range1_w_multipliernode_w_range10569w(0) <= multipliernode_w(54);
	wire_crr_fp_range1_w_multipliernode_w_range10574w(0) <= multipliernode_w(55);
	wire_crr_fp_range1_w_multipliernode_w_range10579w(0) <= multipliernode_w(56);
	wire_crr_fp_range1_w_multipliernode_w_range10584w(0) <= multipliernode_w(57);
	wire_crr_fp_range1_w_multipliernode_w_range10589w(0) <= multipliernode_w(58);
	wire_crr_fp_range1_w_multipliernode_w_range10594w(0) <= multipliernode_w(59);
	wire_crr_fp_range1_w_multipliernode_w_range10324w(0) <= multipliernode_w(5);
	wire_crr_fp_range1_w_multipliernode_w_range10599w(0) <= multipliernode_w(60);
	wire_crr_fp_range1_w_multipliernode_w_range10604w(0) <= multipliernode_w(61);
	wire_crr_fp_range1_w_multipliernode_w_range10609w(0) <= multipliernode_w(62);
	wire_crr_fp_range1_w_multipliernode_w_range10614w(0) <= multipliernode_w(63);
	wire_crr_fp_range1_w_multipliernode_w_range10619w(0) <= multipliernode_w(64);
	wire_crr_fp_range1_w_multipliernode_w_range10624w(0) <= multipliernode_w(65);
	wire_crr_fp_range1_w_multipliernode_w_range10629w(0) <= multipliernode_w(66);
	wire_crr_fp_range1_w_multipliernode_w_range10634w(0) <= multipliernode_w(67);
	wire_crr_fp_range1_w_multipliernode_w_range10639w(0) <= multipliernode_w(68);
	wire_crr_fp_range1_w_multipliernode_w_range10644w(0) <= multipliernode_w(69);
	wire_crr_fp_range1_w_multipliernode_w_range10329w(0) <= multipliernode_w(6);
	wire_crr_fp_range1_w_multipliernode_w_range10649w(0) <= multipliernode_w(70);
	wire_crr_fp_range1_w_multipliernode_w_range10654w(0) <= multipliernode_w(71);
	wire_crr_fp_range1_w_multipliernode_w_range10659w(0) <= multipliernode_w(72);
	wire_crr_fp_range1_w_multipliernode_w_range10664w(0) <= multipliernode_w(73);
	wire_crr_fp_range1_w_multipliernode_w_range10669w(0) <= multipliernode_w(74);
	wire_crr_fp_range1_w_multipliernode_w_range10674w(0) <= multipliernode_w(75);
	wire_crr_fp_range1_w_multipliernode_w_range10679w(0) <= multipliernode_w(76);
	wire_crr_fp_range1_w_multipliernode_w_range10684w(0) <= multipliernode_w(77);
	wire_crr_fp_range1_w_multipliernode_w_range10280w(0) <= multipliernode_w(78);
	wire_crr_fp_range1_w_multipliernode_w_range10334w(0) <= multipliernode_w(7);
	wire_crr_fp_range1_w_multipliernode_w_range10339w(0) <= multipliernode_w(8);
	wire_crr_fp_range1_w_multipliernode_w_range10344w(0) <= multipliernode_w(9);
	fp_range_table1 :  coshw_altfp_sincos_srrt_koa
	  PORT MAP ( 
		address => tableaddressff,
		basefraction => wire_fp_range_table1_basefraction,
		incexponent => wire_fp_range_table1_incexponent,
		incmantissa => wire_fp_range_table1_incmantissa
	  );
	wire_clz23_data <= ( mantissaff & "111111111");
	clz23 :  coshw_altpriority_encoder_qb6
	  PORT MAP ( 
		data => wire_clz23_data,
		q => wire_clz23_q
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN basefractiondelff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN basefractiondelff <= basefractiondelnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN basefractionff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN basefractionff <= basefractionnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_0 <= basefractionff;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_1 <= cbfd_0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_2 <= cbfd_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_3 <= cbfd_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_4 <= cbfd_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN cbfd_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN cbfd_5 <= cbfd_4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN circleff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN circleff <= circlenode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponentff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN exponentff <= wire_crr_fp_range1_w_data_range10272w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN incexponentff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN incexponentff <= incexponentnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN incmantissaff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN incmantissaff <= incmantissanode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN leadff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN leadff <= leadnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissadelff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN mantissadelff <= mantissaff;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissaff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN mantissaff <= wire_crr_fp_range1_w_data_range10271w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissamultiplierff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN mantissamultiplierff <= mantissamultipliernode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN multipliernormff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN multipliernormff <= multipliernormnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN negbasefractiondelff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN negbasefractiondelff <= negbasefractiondelnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN negcircleff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN negcircleff <= negcirclenode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN negrangeexponentff4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN negrangeexponentff4 <= wire_negrangeexponent_sub4_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN negrangeexponentff5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN negrangeexponentff5 <= wire_negrangeexponent_sub5_result;
			END IF;
		END IF;
	END PROCESS;
	loop53 : FOR i IN 0 TO 6 GENERATE 
		wire_negrangeexponentff5_w_lg_w_lg_w_q_range10692w10696w10697w(i) <= wire_negrangeexponentff5_w_lg_w_q_range10692w10696w(0) AND wire_rangeexponentff_5_w_q_range10695w(i);
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 6 GENERATE 
		wire_negrangeexponentff5_w_lg_w_q_range10692w10694w(i) <= wire_negrangeexponentff5_w_q_range10692w(0) AND wire_negrangeexponentff5_w_q_range10693w(i);
	END GENERATE loop54;
	wire_negrangeexponentff5_w_lg_w_q_range10692w10696w(0) <= NOT wire_negrangeexponentff5_w_q_range10692w(0);
	wire_negrangeexponentff5_w_q_range10693w <= negrangeexponentff5(6 DOWNTO 0);
	wire_negrangeexponentff5_w_q_range10692w(0) <= negrangeexponentff5(8);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_0 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_0 <= mantissaexponentnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_1 <= wire_rangeexponent_sub1_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_2 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_2 <= rangeexponentff_1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_3 <= rangeexponentff_2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_4 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_4 <= rangeexponentff_3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rangeexponentff_5 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rangeexponentff_5 <= wire_rangeexponent_sub5_result;
			END IF;
		END IF;
	END PROCESS;
	wire_rangeexponentff_5_w_q_range10695w <= rangeexponentff_5(6 DOWNTO 0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rotateff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rotateff <= rotatenode_w;
			END IF;
		END IF;
	END PROCESS;
	wire_rotateff_w_lg_w_q_range10709w10710w(0) <= NOT wire_rotateff_w_q_range10709w(0);
	wire_rotateff_w_lg_w_q_range10713w10714w(0) <= NOT wire_rotateff_w_q_range10713w(0);
	wire_rotateff_w_lg_w_q_range10716w10717w(0) <= NOT wire_rotateff_w_q_range10716w(0);
	wire_rotateff_w_lg_w_q_range10719w10720w(0) <= NOT wire_rotateff_w_q_range10719w(0);
	wire_rotateff_w_lg_w_q_range10722w10723w(0) <= NOT wire_rotateff_w_q_range10722w(0);
	wire_rotateff_w_lg_w_q_range10725w10726w(0) <= NOT wire_rotateff_w_q_range10725w(0);
	wire_rotateff_w_lg_w_q_range10728w10729w(0) <= NOT wire_rotateff_w_q_range10728w(0);
	wire_rotateff_w_lg_w_q_range10731w10732w(0) <= NOT wire_rotateff_w_q_range10731w(0);
	wire_rotateff_w_lg_w_q_range10734w10735w(0) <= NOT wire_rotateff_w_q_range10734w(0);
	wire_rotateff_w_lg_w_q_range10737w10738w(0) <= NOT wire_rotateff_w_q_range10737w(0);
	wire_rotateff_w_lg_w_q_range10740w10741w(0) <= NOT wire_rotateff_w_q_range10740w(0);
	wire_rotateff_w_lg_w_q_range10743w10744w(0) <= NOT wire_rotateff_w_q_range10743w(0);
	wire_rotateff_w_lg_w_q_range10746w10747w(0) <= NOT wire_rotateff_w_q_range10746w(0);
	wire_rotateff_w_lg_w_q_range10749w10750w(0) <= NOT wire_rotateff_w_q_range10749w(0);
	wire_rotateff_w_lg_w_q_range10752w10753w(0) <= NOT wire_rotateff_w_q_range10752w(0);
	wire_rotateff_w_lg_w_q_range10755w10756w(0) <= NOT wire_rotateff_w_q_range10755w(0);
	wire_rotateff_w_lg_w_q_range10758w10759w(0) <= NOT wire_rotateff_w_q_range10758w(0);
	wire_rotateff_w_lg_w_q_range10761w10762w(0) <= NOT wire_rotateff_w_q_range10761w(0);
	wire_rotateff_w_lg_w_q_range10764w10765w(0) <= NOT wire_rotateff_w_q_range10764w(0);
	wire_rotateff_w_lg_w_q_range10767w10768w(0) <= NOT wire_rotateff_w_q_range10767w(0);
	wire_rotateff_w_lg_w_q_range10770w10771w(0) <= NOT wire_rotateff_w_q_range10770w(0);
	wire_rotateff_w_lg_w_q_range10773w10774w(0) <= NOT wire_rotateff_w_q_range10773w(0);
	wire_rotateff_w_lg_w_q_range10776w10777w(0) <= NOT wire_rotateff_w_q_range10776w(0);
	wire_rotateff_w_lg_w_q_range10779w10780w(0) <= NOT wire_rotateff_w_q_range10779w(0);
	wire_rotateff_w_lg_w_q_range10782w10783w(0) <= NOT wire_rotateff_w_q_range10782w(0);
	wire_rotateff_w_lg_w_q_range10785w10786w(0) <= NOT wire_rotateff_w_q_range10785w(0);
	wire_rotateff_w_lg_w_q_range10788w10789w(0) <= NOT wire_rotateff_w_q_range10788w(0);
	wire_rotateff_w_lg_w_q_range10791w10792w(0) <= NOT wire_rotateff_w_q_range10791w(0);
	wire_rotateff_w_lg_w_q_range10794w10795w(0) <= NOT wire_rotateff_w_q_range10794w(0);
	wire_rotateff_w_lg_w_q_range10797w10798w(0) <= NOT wire_rotateff_w_q_range10797w(0);
	wire_rotateff_w_lg_w_q_range10800w10801w(0) <= NOT wire_rotateff_w_q_range10800w(0);
	wire_rotateff_w_lg_w_q_range10803w10804w(0) <= NOT wire_rotateff_w_q_range10803w(0);
	wire_rotateff_w_lg_w_q_range10806w10807w(0) <= NOT wire_rotateff_w_q_range10806w(0);
	wire_rotateff_w_lg_w_q_range10809w10810w(0) <= NOT wire_rotateff_w_q_range10809w(0);
	wire_rotateff_w_lg_w_q_range10812w10813w(0) <= NOT wire_rotateff_w_q_range10812w(0);
	wire_rotateff_w_lg_w_q_range10815w10816w(0) <= NOT wire_rotateff_w_q_range10815w(0);
	wire_rotateff_w_q_range10709w(0) <= rotateff(42);
	wire_rotateff_w_q_range10713w(0) <= rotateff(43);
	wire_rotateff_w_q_range10716w(0) <= rotateff(44);
	wire_rotateff_w_q_range10719w(0) <= rotateff(45);
	wire_rotateff_w_q_range10722w(0) <= rotateff(46);
	wire_rotateff_w_q_range10725w(0) <= rotateff(47);
	wire_rotateff_w_q_range10728w(0) <= rotateff(48);
	wire_rotateff_w_q_range10731w(0) <= rotateff(49);
	wire_rotateff_w_q_range10734w(0) <= rotateff(50);
	wire_rotateff_w_q_range10737w(0) <= rotateff(51);
	wire_rotateff_w_q_range10740w(0) <= rotateff(52);
	wire_rotateff_w_q_range10743w(0) <= rotateff(53);
	wire_rotateff_w_q_range10746w(0) <= rotateff(54);
	wire_rotateff_w_q_range10749w(0) <= rotateff(55);
	wire_rotateff_w_q_range10752w(0) <= rotateff(56);
	wire_rotateff_w_q_range10755w(0) <= rotateff(57);
	wire_rotateff_w_q_range10758w(0) <= rotateff(58);
	wire_rotateff_w_q_range10761w(0) <= rotateff(59);
	wire_rotateff_w_q_range10764w(0) <= rotateff(60);
	wire_rotateff_w_q_range10767w(0) <= rotateff(61);
	wire_rotateff_w_q_range10770w(0) <= rotateff(62);
	wire_rotateff_w_q_range10773w(0) <= rotateff(63);
	wire_rotateff_w_q_range10776w(0) <= rotateff(64);
	wire_rotateff_w_q_range10779w(0) <= rotateff(65);
	wire_rotateff_w_q_range10782w(0) <= rotateff(66);
	wire_rotateff_w_q_range10785w(0) <= rotateff(67);
	wire_rotateff_w_q_range10788w(0) <= rotateff(68);
	wire_rotateff_w_q_range10791w(0) <= rotateff(69);
	wire_rotateff_w_q_range10794w(0) <= rotateff(70);
	wire_rotateff_w_q_range10797w(0) <= rotateff(71);
	wire_rotateff_w_q_range10800w(0) <= rotateff(72);
	wire_rotateff_w_q_range10803w(0) <= rotateff(73);
	wire_rotateff_w_q_range10806w(0) <= rotateff(74);
	wire_rotateff_w_q_range10809w(0) <= rotateff(75);
	wire_rotateff_w_q_range10812w(0) <= rotateff(76);
	wire_rotateff_w_q_range10815w(0) <= rotateff(77);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN tableaddressff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN tableaddressff <= exponentff;
			END IF;
		END IF;
	END PROCESS;
	wire_circle_add_dataa <= ( "0" & basefractiondelff);
	wire_circle_add_datab <= ( "0" & rotateff(77 DOWNTO 42));
	circle_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 37
	  )
	  PORT MAP ( 
		dataa => wire_circle_add_dataa,
		datab => wire_circle_add_datab,
		result => wire_circle_add_result
	  );
	wire_exponent_adjust_sub_datab <= ( "0000" & leadff);
	exponent_adjust_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => const_23_w,
		datab => wire_exponent_adjust_sub_datab,
		result => wire_exponent_adjust_sub_result
	  );
	wire_negbasedractiondel_sub_dataa <= (OTHERS => '0');
	negbasedractiondel_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 36
	  )
	  PORT MAP ( 
		dataa => wire_negbasedractiondel_sub_dataa,
		datab => basefractiondelnode_w(35 DOWNTO 0),
		result => wire_negbasedractiondel_sub_result
	  );
	wire_negcircle_add_dataa <= ( "1" & negbasefractiondelff);
	wire_negcircle_add_datab <= ( "1" & negrotatenode_w);
	negcircle_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 37
	  )
	  PORT MAP ( 
		cin => wire_vcc,
		dataa => wire_negcircle_add_dataa,
		datab => wire_negcircle_add_datab,
		result => wire_negcircle_add_result
	  );
	wire_negrangeexponent_sub4_dataa <= ( "1" & "00000000");
	negrangeexponent_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => wire_negrangeexponent_sub4_dataa,
		datab => rangeexponentff_3,
		result => wire_negrangeexponent_sub4_result
	  );
	wire_negrangeexponent_sub5_datab <= ( "00000000" & wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w);
	negrangeexponent_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => negrangeexponentff4,
		datab => wire_negrangeexponent_sub5_datab,
		result => wire_negrangeexponent_sub5_result
	  );
	wire_rangeexponent_sub1_datab <= ( "0" & incexponentff);
	rangeexponent_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => rangeexponentff_0,
		datab => wire_rangeexponent_sub1_datab,
		result => wire_rangeexponent_sub1_result
	  );
	wire_rangeexponent_sub5_datab <= ( "00000000" & wire_crr_fp_range1_w_lg_w_multipliernode_w_range10280w10281w);
	rangeexponent_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => rangeexponentff_4,
		datab => wire_rangeexponent_sub5_datab,
		result => wire_rangeexponent_sub5_result
	  );
	csftin :  lpm_clshift
	  GENERIC MAP (
		LPM_WIDTH => 23,
		LPM_WIDTHDIST => 5
	  )
	  PORT MAP ( 
		data => mantissadelff,
		direction => wire_gnd,
		distance => leadff,
		result => wire_csftin_result
	  );
	wire_fp_lsft_rsft78_distance <= wire_negrangeexponentff5_w_lg_w_lg_w_lg_w_q_range10692w10696w10697w10698w;
	loop55 : FOR i IN 0 TO 6 GENERATE 
		wire_negrangeexponentff5_w_lg_w_lg_w_lg_w_q_range10692w10696w10697w10698w(i) <= wire_negrangeexponentff5_w_lg_w_lg_w_q_range10692w10696w10697w(i) OR wire_negrangeexponentff5_w_lg_w_q_range10692w10694w(i);
	END GENERATE loop55;
	fp_lsft_rsft78 :  lpm_clshift
	  GENERIC MAP (
		LPM_PIPELINE => 1,
		LPM_WIDTH => 78,
		LPM_WIDTHDIST => 7
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		data => multipliernormff,
		direction => negrangeexponentff5(8),
		distance => wire_fp_lsft_rsft78_distance,
		result => wire_fp_lsft_rsft78_result
	  );
	mult23x56 :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 4,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 23,
		LPM_WIDTHB => 56,
		LPM_WIDTHP => 79
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => mantissamultiplierff,
		datab => incmantissaff,
		result => wire_mult23x56_result
	  );

 END RTL; --coshw_altfp_sincos_range_b6c


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" WIDTH=64 WIDTHAD=6 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=32 WIDTHAD=5 data q
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altpriority_encoder_q08 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0)
	 ); 
 END coshw_altpriority_encoder_q08;

 ARCHITECTURE RTL OF coshw_altpriority_encoder_q08 IS

	 SIGNAL  wire_altpriority_encoder19_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero12306w12307w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero12308w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_zero12306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_w_lg_w_lg_zero12308w12309w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder20_zero	:	STD_LOGIC;
	 COMPONENT  coshw_altpriority_encoder_r08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder20_w_lg_zero12306w & wire_altpriority_encoder20_w_lg_w_lg_zero12308w12309w);
	altpriority_encoder19 :  coshw_altpriority_encoder_r08
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder19_q
	  );
	loop56 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero12306w12307w(i) <= wire_altpriority_encoder20_w_lg_zero12306w(0) AND wire_altpriority_encoder20_q(i);
	END GENERATE loop56;
	loop57 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder20_w_lg_zero12308w(i) <= wire_altpriority_encoder20_zero AND wire_altpriority_encoder19_q(i);
	END GENERATE loop57;
	wire_altpriority_encoder20_w_lg_zero12306w(0) <= NOT wire_altpriority_encoder20_zero;
	loop58 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder20_w_lg_w_lg_zero12308w12309w(i) <= wire_altpriority_encoder20_w_lg_zero12308w(i) OR wire_altpriority_encoder20_w_lg_w_lg_zero12306w12307w(i);
	END GENERATE loop58;
	altpriority_encoder20 :  coshw_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder20_q,
		zero => wire_altpriority_encoder20_zero
	  );

 END RTL; --coshw_altpriority_encoder_q08


--altpriority_encoder CBX_AUTO_BLACKBOX="ALL" LSB_PRIORITY="NO" WIDTH=32 WIDTHAD=5 data q zero
--VERSION_BEGIN 18.1 cbx_altpriority_encoder 2018:09:12:13:04:24:SJ cbx_mgl 2018:09:12:13:10:36:SJ  VERSION_END

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altpriority_encoder_qf8 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 zero	:	OUT  STD_LOGIC
	 ); 
 END coshw_altpriority_encoder_qf8;

 ARCHITECTURE RTL OF coshw_altpriority_encoder_qf8 IS

	 SIGNAL  wire_altpriority_encoder21_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder21_zero	:	STD_LOGIC;
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero12315w12316w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero12317w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_zero12315w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_w_lg_w_lg_zero12317w12318w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_q	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder22_zero	:	STD_LOGIC;
	 COMPONENT  coshw_altpriority_encoder_rf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(3 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder22_w_lg_zero12315w & wire_altpriority_encoder22_w_lg_w_lg_zero12317w12318w);
	zero <= (wire_altpriority_encoder21_zero AND wire_altpriority_encoder22_zero);
	altpriority_encoder21 :  coshw_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(15 DOWNTO 0),
		q => wire_altpriority_encoder21_q,
		zero => wire_altpriority_encoder21_zero
	  );
	loop59 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder22_w_lg_w_lg_zero12315w12316w(i) <= wire_altpriority_encoder22_w_lg_zero12315w(0) AND wire_altpriority_encoder22_q(i);
	END GENERATE loop59;
	loop60 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder22_w_lg_zero12317w(i) <= wire_altpriority_encoder22_zero AND wire_altpriority_encoder21_q(i);
	END GENERATE loop60;
	wire_altpriority_encoder22_w_lg_zero12315w(0) <= NOT wire_altpriority_encoder22_zero;
	loop61 : FOR i IN 0 TO 3 GENERATE 
		wire_altpriority_encoder22_w_lg_w_lg_zero12317w12318w(i) <= wire_altpriority_encoder22_w_lg_zero12317w(i) OR wire_altpriority_encoder22_w_lg_w_lg_zero12315w12316w(i);
	END GENERATE loop61;
	altpriority_encoder22 :  coshw_altpriority_encoder_rf8
	  PORT MAP ( 
		data => data(31 DOWNTO 16),
		q => wire_altpriority_encoder22_q,
		zero => wire_altpriority_encoder22_zero
	  );

 END RTL; --coshw_altpriority_encoder_qf8

--synthesis_resources = 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altpriority_encoder_0c6 IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 q	:	OUT  STD_LOGIC_VECTOR (5 DOWNTO 0)
	 ); 
 END coshw_altpriority_encoder_0c6;

 ARCHITECTURE RTL OF coshw_altpriority_encoder_0c6 IS

	 SIGNAL  wire_altpriority_encoder17_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero12297w12298w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero12299w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_zero12297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_w_lg_w_lg_zero12299w12300w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_q	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_altpriority_encoder18_zero	:	STD_LOGIC;
	 COMPONENT  coshw_altpriority_encoder_q08
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altpriority_encoder_qf8
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(4 DOWNTO 0);
		zero	:	OUT  STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	q <= ( wire_altpriority_encoder18_w_lg_zero12297w & wire_altpriority_encoder18_w_lg_w_lg_zero12299w12300w);
	altpriority_encoder17 :  coshw_altpriority_encoder_q08
	  PORT MAP ( 
		data => data(31 DOWNTO 0),
		q => wire_altpriority_encoder17_q
	  );
	loop62 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder18_w_lg_w_lg_zero12297w12298w(i) <= wire_altpriority_encoder18_w_lg_zero12297w(0) AND wire_altpriority_encoder18_q(i);
	END GENERATE loop62;
	loop63 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder18_w_lg_zero12299w(i) <= wire_altpriority_encoder18_zero AND wire_altpriority_encoder17_q(i);
	END GENERATE loop63;
	wire_altpriority_encoder18_w_lg_zero12297w(0) <= NOT wire_altpriority_encoder18_zero;
	loop64 : FOR i IN 0 TO 4 GENERATE 
		wire_altpriority_encoder18_w_lg_w_lg_zero12299w12300w(i) <= wire_altpriority_encoder18_w_lg_zero12299w(i) OR wire_altpriority_encoder18_w_lg_w_lg_zero12297w12298w(i);
	END GENERATE loop64;
	altpriority_encoder18 :  coshw_altpriority_encoder_qf8
	  PORT MAP ( 
		data => data(63 DOWNTO 32),
		q => wire_altpriority_encoder18_q,
		zero => wire_altpriority_encoder18_zero
	  );

 END RTL; --coshw_altpriority_encoder_0c6

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 51 lpm_clshift 3 lpm_mult 3 lpm_mux 2 reg 2434 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  coshw_altfp_sincos_u6e IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 data	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END coshw_altfp_sincos_u6e;

 ARCHITECTURE RTL OF coshw_altfp_sincos_u6e IS

	 SIGNAL  wire_ccc_cordic_m_sincos	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_circle	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_crr_fp_range1_negcircle	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_clz_data	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_clz_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL	 countff	:	STD_LOGIC_VECTOR(5 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exponentnormff	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 fixed_sincosff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 mantissanormff	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 quadrant_sumff	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 select_sincosff	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 signcalcff	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 signinff	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exponentnorm_add_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exponentnorm_add_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exponentnormmode_sub_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_exponentnormmode_sub_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_mantissanorm_add_datab	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_mantissanorm_add_result	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_quadrantsum_add_result	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_sft_result	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_cmul_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_negative_quadrant_w23w	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_w_lg_positive_quadrant_w24w	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_circle_w_range11w12w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_circle_w_range3w4w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range204w205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range207w208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range210w211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range213w214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range216w217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range219w220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range222w223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range225w226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range228w229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range231w232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range234w235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range237w238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range240w241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range243w244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range246w247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range249w250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range252w253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range255w256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range258w259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range261w262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range264w265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range267w268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_mantissanormnode_w_range270w271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_negcircle_w_range8w9w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_lg_quadrantselect_w10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_circle_w_range1w2w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_quadrant_w_range21w22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range142w144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range172w174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range175w177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range178w180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range181w183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range184w186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range145w147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range148w150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range151w153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range154w156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range157w159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range160w162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range163w165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range166w168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_indexcheck_w_range169w171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  circle_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  countnode_w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  exponentnormmode_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  fixed_sincos_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  fixed_sincosnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  fraction_quadrant_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  indexbit_w :	STD_LOGIC;
	 SIGNAL  indexcheck_w :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  mantissanormnode_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  negative_quadrant_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  negcircle_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  one_term_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  overflownode_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  piovertwo_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  positive_quadrant_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  quadrant_w :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  quadrantselect_w :	STD_LOGIC;
	 SIGNAL  quadrantsign_w :	STD_LOGIC;
	 SIGNAL  radiansnode_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  value_128_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  zerovec_w :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_w_circle_w_range11w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_circle_w_range1w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_circle_w_range3w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_indexcheck_w_range169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_mantissanormnode_w_range270w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_negcircle_w_range8w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_overflownode_w_range230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_quadrant_w_range21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_radiansnode_w_range141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  coshw_altfp_sincos_cordic_m_d5e
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		indexbit	:	IN  STD_LOGIC := '0';
		radians	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
		sincos	:	OUT  STD_LOGIC_VECTOR(31 DOWNTO 0);
		sincosbit	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altfp_sincos_range_b6c
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		circle	:	OUT  STD_LOGIC_VECTOR(35 DOWNTO 0);
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		data	:	IN  STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
		negcircle	:	OUT  STD_LOGIC_VECTOR(35 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  coshw_altpriority_encoder_0c6
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(63 DOWNTO 0);
		q	:	OUT  STD_LOGIC_VECTOR(5 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_clshift
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_SHIFTTYPE	:	STRING := "LOGICAL";
		LPM_WIDTH	:	NATURAL;
		LPM_WIDTHDIST	:	NATURAL;
		lpm_type	:	STRING := "lpm_clshift"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		direction	:	IN STD_LOGIC := '0';
		distance	:	IN STD_LOGIC_VECTOR(LPM_WIDTHDIST-1 DOWNTO 0);
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		underflow	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_mult
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTHA	:	NATURAL;
		LPM_WIDTHB	:	NATURAL;
		LPM_WIDTHP	:	NATURAL;
		LPM_WIDTHS	:	NATURAL := 1;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_mult"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTHA-1 DOWNTO 0);
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTHB-1 DOWNTO 0);
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTHP-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sum	:	IN STD_LOGIC_VECTOR(LPM_WIDTHS-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	loop65 : FOR i IN 0 TO 35 GENERATE 
		wire_w_lg_negative_quadrant_w23w(i) <= negative_quadrant_w(i) AND wire_w_lg_w_quadrant_w_range21w22w(0);
	END GENERATE loop65;
	loop66 : FOR i IN 0 TO 35 GENERATE 
		wire_w_lg_positive_quadrant_w24w(i) <= positive_quadrant_w(i) AND wire_w_quadrant_w_range21w(0);
	END GENERATE loop66;
	loop67 : FOR i IN 0 TO 33 GENERATE 
		wire_w_lg_w_circle_w_range11w12w(i) <= wire_w_circle_w_range11w(i) AND wire_w_lg_quadrantselect_w10w(0);
	END GENERATE loop67;
	wire_w_lg_w_circle_w_range3w4w(0) <= wire_w_circle_w_range3w(0) AND wire_w_lg_w_circle_w_range1w2w(0);
	wire_w_lg_w_mantissanormnode_w_range204w205w(0) <= wire_w_mantissanormnode_w_range204w(0) AND wire_w_overflownode_w_range202w(0);
	wire_w_lg_w_mantissanormnode_w_range207w208w(0) <= wire_w_mantissanormnode_w_range207w(0) AND wire_w_overflownode_w_range206w(0);
	wire_w_lg_w_mantissanormnode_w_range210w211w(0) <= wire_w_mantissanormnode_w_range210w(0) AND wire_w_overflownode_w_range209w(0);
	wire_w_lg_w_mantissanormnode_w_range213w214w(0) <= wire_w_mantissanormnode_w_range213w(0) AND wire_w_overflownode_w_range212w(0);
	wire_w_lg_w_mantissanormnode_w_range216w217w(0) <= wire_w_mantissanormnode_w_range216w(0) AND wire_w_overflownode_w_range215w(0);
	wire_w_lg_w_mantissanormnode_w_range219w220w(0) <= wire_w_mantissanormnode_w_range219w(0) AND wire_w_overflownode_w_range218w(0);
	wire_w_lg_w_mantissanormnode_w_range222w223w(0) <= wire_w_mantissanormnode_w_range222w(0) AND wire_w_overflownode_w_range221w(0);
	wire_w_lg_w_mantissanormnode_w_range225w226w(0) <= wire_w_mantissanormnode_w_range225w(0) AND wire_w_overflownode_w_range224w(0);
	wire_w_lg_w_mantissanormnode_w_range228w229w(0) <= wire_w_mantissanormnode_w_range228w(0) AND wire_w_overflownode_w_range227w(0);
	wire_w_lg_w_mantissanormnode_w_range231w232w(0) <= wire_w_mantissanormnode_w_range231w(0) AND wire_w_overflownode_w_range230w(0);
	wire_w_lg_w_mantissanormnode_w_range234w235w(0) <= wire_w_mantissanormnode_w_range234w(0) AND wire_w_overflownode_w_range233w(0);
	wire_w_lg_w_mantissanormnode_w_range237w238w(0) <= wire_w_mantissanormnode_w_range237w(0) AND wire_w_overflownode_w_range236w(0);
	wire_w_lg_w_mantissanormnode_w_range240w241w(0) <= wire_w_mantissanormnode_w_range240w(0) AND wire_w_overflownode_w_range239w(0);
	wire_w_lg_w_mantissanormnode_w_range243w244w(0) <= wire_w_mantissanormnode_w_range243w(0) AND wire_w_overflownode_w_range242w(0);
	wire_w_lg_w_mantissanormnode_w_range246w247w(0) <= wire_w_mantissanormnode_w_range246w(0) AND wire_w_overflownode_w_range245w(0);
	wire_w_lg_w_mantissanormnode_w_range249w250w(0) <= wire_w_mantissanormnode_w_range249w(0) AND wire_w_overflownode_w_range248w(0);
	wire_w_lg_w_mantissanormnode_w_range252w253w(0) <= wire_w_mantissanormnode_w_range252w(0) AND wire_w_overflownode_w_range251w(0);
	wire_w_lg_w_mantissanormnode_w_range255w256w(0) <= wire_w_mantissanormnode_w_range255w(0) AND wire_w_overflownode_w_range254w(0);
	wire_w_lg_w_mantissanormnode_w_range258w259w(0) <= wire_w_mantissanormnode_w_range258w(0) AND wire_w_overflownode_w_range257w(0);
	wire_w_lg_w_mantissanormnode_w_range261w262w(0) <= wire_w_mantissanormnode_w_range261w(0) AND wire_w_overflownode_w_range260w(0);
	wire_w_lg_w_mantissanormnode_w_range264w265w(0) <= wire_w_mantissanormnode_w_range264w(0) AND wire_w_overflownode_w_range263w(0);
	wire_w_lg_w_mantissanormnode_w_range267w268w(0) <= wire_w_mantissanormnode_w_range267w(0) AND wire_w_overflownode_w_range266w(0);
	wire_w_lg_w_mantissanormnode_w_range270w271w(0) <= wire_w_mantissanormnode_w_range270w(0) AND wire_w_overflownode_w_range269w(0);
	loop68 : FOR i IN 0 TO 33 GENERATE 
		wire_w_lg_w_negcircle_w_range8w9w(i) <= wire_w_negcircle_w_range8w(i) AND quadrantselect_w;
	END GENERATE loop68;
	wire_w_lg_quadrantselect_w10w(0) <= NOT quadrantselect_w;
	wire_w_lg_w_circle_w_range1w2w(0) <= NOT wire_w_circle_w_range1w(0);
	wire_w_lg_w_quadrant_w_range21w22w(0) <= NOT wire_w_quadrant_w_range21w(0);
	wire_w_lg_w_indexcheck_w_range142w144w(0) <= wire_w_indexcheck_w_range142w(0) OR wire_w_radiansnode_w_range141w(0);
	wire_w_lg_w_indexcheck_w_range172w174w(0) <= wire_w_indexcheck_w_range172w(0) OR wire_w_radiansnode_w_range173w(0);
	wire_w_lg_w_indexcheck_w_range175w177w(0) <= wire_w_indexcheck_w_range175w(0) OR wire_w_radiansnode_w_range176w(0);
	wire_w_lg_w_indexcheck_w_range178w180w(0) <= wire_w_indexcheck_w_range178w(0) OR wire_w_radiansnode_w_range179w(0);
	wire_w_lg_w_indexcheck_w_range181w183w(0) <= wire_w_indexcheck_w_range181w(0) OR wire_w_radiansnode_w_range182w(0);
	wire_w_lg_w_indexcheck_w_range184w186w(0) <= wire_w_indexcheck_w_range184w(0) OR wire_w_radiansnode_w_range185w(0);
	wire_w_lg_w_indexcheck_w_range145w147w(0) <= wire_w_indexcheck_w_range145w(0) OR wire_w_radiansnode_w_range146w(0);
	wire_w_lg_w_indexcheck_w_range148w150w(0) <= wire_w_indexcheck_w_range148w(0) OR wire_w_radiansnode_w_range149w(0);
	wire_w_lg_w_indexcheck_w_range151w153w(0) <= wire_w_indexcheck_w_range151w(0) OR wire_w_radiansnode_w_range152w(0);
	wire_w_lg_w_indexcheck_w_range154w156w(0) <= wire_w_indexcheck_w_range154w(0) OR wire_w_radiansnode_w_range155w(0);
	wire_w_lg_w_indexcheck_w_range157w159w(0) <= wire_w_indexcheck_w_range157w(0) OR wire_w_radiansnode_w_range158w(0);
	wire_w_lg_w_indexcheck_w_range160w162w(0) <= wire_w_indexcheck_w_range160w(0) OR wire_w_radiansnode_w_range161w(0);
	wire_w_lg_w_indexcheck_w_range163w165w(0) <= wire_w_indexcheck_w_range163w(0) OR wire_w_radiansnode_w_range164w(0);
	wire_w_lg_w_indexcheck_w_range166w168w(0) <= wire_w_indexcheck_w_range166w(0) OR wire_w_radiansnode_w_range167w(0);
	wire_w_lg_w_indexcheck_w_range169w171w(0) <= wire_w_indexcheck_w_range169w(0) OR wire_w_radiansnode_w_range170w(0);
	aclr <= '0';
	circle_w <= wire_crr_fp_range1_circle;
	clk_en <= '1';
	countnode_w <= (NOT wire_clz_q);
	exponentnormmode_w <= wire_exponentnormmode_sub_result;
	fixed_sincos_w <= wire_ccc_cordic_m_sincos;
	fixed_sincosnode_w <= ( fixed_sincos_w & zerovec_w(3 DOWNTO 0));
	fraction_quadrant_w <= (wire_w_lg_positive_quadrant_w24w OR wire_w_lg_negative_quadrant_w23w);
	indexbit_w <= (NOT indexcheck_w(4));
	indexcheck_w <= ( wire_w_lg_w_indexcheck_w_range184w186w & wire_w_lg_w_indexcheck_w_range181w183w & wire_w_lg_w_indexcheck_w_range178w180w & wire_w_lg_w_indexcheck_w_range175w177w & wire_w_lg_w_indexcheck_w_range172w174w & wire_w_lg_w_indexcheck_w_range169w171w & wire_w_lg_w_indexcheck_w_range166w168w & wire_w_lg_w_indexcheck_w_range163w165w & wire_w_lg_w_indexcheck_w_range160w162w & wire_w_lg_w_indexcheck_w_range157w159w & wire_w_lg_w_indexcheck_w_range154w156w & wire_w_lg_w_indexcheck_w_range151w153w & wire_w_lg_w_indexcheck_w_range148w150w & wire_w_lg_w_indexcheck_w_range145w147w & wire_w_lg_w_indexcheck_w_range142w144w & radiansnode_w(30));
	mantissanormnode_w <= wire_sft_result;
	negative_quadrant_w <= (NOT positive_quadrant_w);
	negcircle_w <= wire_crr_fp_range1_negcircle;
	one_term_w <= ( wire_w_lg_w_quadrant_w_range21w22w & zerovec_w(34 DOWNTO 0));
	overflownode_w <= ( wire_w_lg_w_mantissanormnode_w_range270w271w & wire_w_lg_w_mantissanormnode_w_range267w268w & wire_w_lg_w_mantissanormnode_w_range264w265w & wire_w_lg_w_mantissanormnode_w_range261w262w & wire_w_lg_w_mantissanormnode_w_range258w259w & wire_w_lg_w_mantissanormnode_w_range255w256w & wire_w_lg_w_mantissanormnode_w_range252w253w & wire_w_lg_w_mantissanormnode_w_range249w250w & wire_w_lg_w_mantissanormnode_w_range246w247w & wire_w_lg_w_mantissanormnode_w_range243w244w & wire_w_lg_w_mantissanormnode_w_range240w241w & wire_w_lg_w_mantissanormnode_w_range237w238w & wire_w_lg_w_mantissanormnode_w_range234w235w & wire_w_lg_w_mantissanormnode_w_range231w232w & wire_w_lg_w_mantissanormnode_w_range228w229w & wire_w_lg_w_mantissanormnode_w_range225w226w & wire_w_lg_w_mantissanormnode_w_range222w223w & wire_w_lg_w_mantissanormnode_w_range219w220w & wire_w_lg_w_mantissanormnode_w_range216w217w & wire_w_lg_w_mantissanormnode_w_range213w214w & wire_w_lg_w_mantissanormnode_w_range210w211w & wire_w_lg_w_mantissanormnode_w_range207w208w & wire_w_lg_w_mantissanormnode_w_range204w205w & mantissanormnode_w(11));
	piovertwo_w <= "110010010000111111011010101000100010";
	positive_quadrant_w <= ( "0" & quadrant_w & "0");
	quadrant_w <= (wire_w_lg_w_circle_w_range11w12w OR wire_w_lg_w_negcircle_w_range8w9w);
	quadrantselect_w <= circle_w(34);
	quadrantsign_w <= (((NOT circle_w(35)) AND circle_w(34)) OR wire_w_lg_w_circle_w_range3w4w(0));
	radiansnode_w <= wire_cmul_result;
	result <= ( signcalcff(23) & exponentnormff & mantissanormff);
	value_128_w <= "10000000";
	zerovec_w <= (OTHERS => '0');
	wire_w_circle_w_range11w <= circle_w(33 DOWNTO 0);
	wire_w_circle_w_range1w(0) <= circle_w(34);
	wire_w_circle_w_range3w(0) <= circle_w(35);
	wire_w_indexcheck_w_range142w(0) <= indexcheck_w(0);
	wire_w_indexcheck_w_range172w(0) <= indexcheck_w(10);
	wire_w_indexcheck_w_range175w(0) <= indexcheck_w(11);
	wire_w_indexcheck_w_range178w(0) <= indexcheck_w(12);
	wire_w_indexcheck_w_range181w(0) <= indexcheck_w(13);
	wire_w_indexcheck_w_range184w(0) <= indexcheck_w(14);
	wire_w_indexcheck_w_range145w(0) <= indexcheck_w(1);
	wire_w_indexcheck_w_range148w(0) <= indexcheck_w(2);
	wire_w_indexcheck_w_range151w(0) <= indexcheck_w(3);
	wire_w_indexcheck_w_range154w(0) <= indexcheck_w(4);
	wire_w_indexcheck_w_range157w(0) <= indexcheck_w(5);
	wire_w_indexcheck_w_range160w(0) <= indexcheck_w(6);
	wire_w_indexcheck_w_range163w(0) <= indexcheck_w(7);
	wire_w_indexcheck_w_range166w(0) <= indexcheck_w(8);
	wire_w_indexcheck_w_range169w(0) <= indexcheck_w(9);
	wire_w_mantissanormnode_w_range204w(0) <= mantissanormnode_w(12);
	wire_w_mantissanormnode_w_range207w(0) <= mantissanormnode_w(13);
	wire_w_mantissanormnode_w_range210w(0) <= mantissanormnode_w(14);
	wire_w_mantissanormnode_w_range213w(0) <= mantissanormnode_w(15);
	wire_w_mantissanormnode_w_range216w(0) <= mantissanormnode_w(16);
	wire_w_mantissanormnode_w_range219w(0) <= mantissanormnode_w(17);
	wire_w_mantissanormnode_w_range222w(0) <= mantissanormnode_w(18);
	wire_w_mantissanormnode_w_range225w(0) <= mantissanormnode_w(19);
	wire_w_mantissanormnode_w_range228w(0) <= mantissanormnode_w(20);
	wire_w_mantissanormnode_w_range231w(0) <= mantissanormnode_w(21);
	wire_w_mantissanormnode_w_range234w(0) <= mantissanormnode_w(22);
	wire_w_mantissanormnode_w_range237w(0) <= mantissanormnode_w(23);
	wire_w_mantissanormnode_w_range240w(0) <= mantissanormnode_w(24);
	wire_w_mantissanormnode_w_range243w(0) <= mantissanormnode_w(25);
	wire_w_mantissanormnode_w_range246w(0) <= mantissanormnode_w(26);
	wire_w_mantissanormnode_w_range249w(0) <= mantissanormnode_w(27);
	wire_w_mantissanormnode_w_range252w(0) <= mantissanormnode_w(28);
	wire_w_mantissanormnode_w_range255w(0) <= mantissanormnode_w(29);
	wire_w_mantissanormnode_w_range258w(0) <= mantissanormnode_w(30);
	wire_w_mantissanormnode_w_range261w(0) <= mantissanormnode_w(31);
	wire_w_mantissanormnode_w_range264w(0) <= mantissanormnode_w(32);
	wire_w_mantissanormnode_w_range267w(0) <= mantissanormnode_w(33);
	wire_w_mantissanormnode_w_range270w(0) <= mantissanormnode_w(34);
	wire_w_negcircle_w_range8w <= negcircle_w(33 DOWNTO 0);
	wire_w_overflownode_w_range202w(0) <= overflownode_w(0);
	wire_w_overflownode_w_range233w(0) <= overflownode_w(10);
	wire_w_overflownode_w_range236w(0) <= overflownode_w(11);
	wire_w_overflownode_w_range239w(0) <= overflownode_w(12);
	wire_w_overflownode_w_range242w(0) <= overflownode_w(13);
	wire_w_overflownode_w_range245w(0) <= overflownode_w(14);
	wire_w_overflownode_w_range248w(0) <= overflownode_w(15);
	wire_w_overflownode_w_range251w(0) <= overflownode_w(16);
	wire_w_overflownode_w_range254w(0) <= overflownode_w(17);
	wire_w_overflownode_w_range257w(0) <= overflownode_w(18);
	wire_w_overflownode_w_range260w(0) <= overflownode_w(19);
	wire_w_overflownode_w_range206w(0) <= overflownode_w(1);
	wire_w_overflownode_w_range263w(0) <= overflownode_w(20);
	wire_w_overflownode_w_range266w(0) <= overflownode_w(21);
	wire_w_overflownode_w_range269w(0) <= overflownode_w(22);
	wire_w_overflownode_w_range209w(0) <= overflownode_w(2);
	wire_w_overflownode_w_range212w(0) <= overflownode_w(3);
	wire_w_overflownode_w_range215w(0) <= overflownode_w(4);
	wire_w_overflownode_w_range218w(0) <= overflownode_w(5);
	wire_w_overflownode_w_range221w(0) <= overflownode_w(6);
	wire_w_overflownode_w_range224w(0) <= overflownode_w(7);
	wire_w_overflownode_w_range227w(0) <= overflownode_w(8);
	wire_w_overflownode_w_range230w(0) <= overflownode_w(9);
	wire_w_quadrant_w_range21w(0) <= quadrant_w(33);
	wire_w_radiansnode_w_range185w(0) <= radiansnode_w(16);
	wire_w_radiansnode_w_range182w(0) <= radiansnode_w(17);
	wire_w_radiansnode_w_range179w(0) <= radiansnode_w(18);
	wire_w_radiansnode_w_range176w(0) <= radiansnode_w(19);
	wire_w_radiansnode_w_range173w(0) <= radiansnode_w(20);
	wire_w_radiansnode_w_range170w(0) <= radiansnode_w(21);
	wire_w_radiansnode_w_range167w(0) <= radiansnode_w(22);
	wire_w_radiansnode_w_range164w(0) <= radiansnode_w(23);
	wire_w_radiansnode_w_range161w(0) <= radiansnode_w(24);
	wire_w_radiansnode_w_range158w(0) <= radiansnode_w(25);
	wire_w_radiansnode_w_range155w(0) <= radiansnode_w(26);
	wire_w_radiansnode_w_range152w(0) <= radiansnode_w(27);
	wire_w_radiansnode_w_range149w(0) <= radiansnode_w(28);
	wire_w_radiansnode_w_range146w(0) <= radiansnode_w(29);
	wire_w_radiansnode_w_range141w(0) <= radiansnode_w(30);
	ccc_cordic_m :  coshw_altfp_sincos_cordic_m_d5e
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		indexbit => indexbit_w,
		radians => radiansnode_w,
		sincos => wire_ccc_cordic_m_sincos,
		sincosbit => select_sincosff(3)
	  );
	crr_fp_range1 :  coshw_altfp_sincos_range_b6c
	  PORT MAP ( 
		aclr => aclr,
		circle => wire_crr_fp_range1_circle,
		clken => clk_en,
		clock => clock,
		data => data,
		negcircle => wire_crr_fp_range1_negcircle
	  );
	wire_clz_data <= ( fixed_sincosnode_w & "1111111111111111111111111111");
	clz :  coshw_altpriority_encoder_0c6
	  PORT MAP ( 
		data => wire_clz_data,
		q => wire_clz_q
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN countff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN countff <= countnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exponentnormff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exponentnormff <= wire_exponentnorm_add_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN fixed_sincosff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN fixed_sincosff <= fixed_sincosnode_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN mantissanormff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN mantissanormff <= wire_mantissanorm_add_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN quadrant_sumff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN quadrant_sumff <= wire_quadrantsum_add_result;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN select_sincosff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN select_sincosff <= ( select_sincosff(2 DOWNTO 0) & wire_w_lg_w_quadrant_w_range21w22w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN signcalcff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN signcalcff <= ( signcalcff(22 DOWNTO 0) & quadrantsign_w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN signinff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN signinff <= ( signinff(9 DOWNTO 0) & data(31));
			END IF;
		END IF;
	END PROCESS;
	wire_exponentnorm_add_datab <= ( "0000000" & overflownode_w(23));
	exponentnorm_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		dataa => exponentnormmode_w(7 DOWNTO 0),
		datab => wire_exponentnorm_add_datab,
		result => wire_exponentnorm_add_result
	  );
	wire_exponentnormmode_sub_datab <= ( "00" & countff);
	exponentnormmode_sub :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		dataa => value_128_w,
		datab => wire_exponentnormmode_sub_datab,
		result => wire_exponentnormmode_sub_result
	  );
	wire_mantissanorm_add_datab <= ( "0000000000000000000000" & mantissanormnode_w(11));
	mantissanorm_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 23
	  )
	  PORT MAP ( 
		dataa => mantissanormnode_w(34 DOWNTO 12),
		datab => wire_mantissanorm_add_datab,
		result => wire_mantissanorm_add_result
	  );
	quadrantsum_add :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 36
	  )
	  PORT MAP ( 
		cin => quadrant_w(33),
		dataa => one_term_w,
		datab => fraction_quadrant_w,
		result => wire_quadrantsum_add_result
	  );
	sft :  lpm_clshift
	  GENERIC MAP (
		LPM_WIDTH => 36,
		LPM_WIDTHDIST => 6
	  )
	  PORT MAP ( 
		data => fixed_sincosff,
		direction => wire_gnd,
		distance => countff,
		result => wire_sft_result
	  );
	cmul :  lpm_mult
	  GENERIC MAP (
		LPM_PIPELINE => 3,
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTHA => 36,
		LPM_WIDTHB => 36,
		LPM_WIDTHP => 32
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => quadrant_sumff,
		datab => piovertwo_w,
		result => wire_cmul_result
	  );

 END RTL; --coshw_altfp_sincos_u6e
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY coshw IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END coshw;


ARCHITECTURE RTL OF coshw IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT coshw_altfp_sincos_u6e
	PORT (
			clock	: IN STD_LOGIC ;
			data	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(31 DOWNTO 0);

	coshw_altfp_sincos_u6e_component : coshw_altfp_sincos_u6e
	PORT MAP (
		clock => clock,
		data => data,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: FPM_FORMAT NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
-- Retrieval info: CONSTANT: OPERATION STRING "COS"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "35"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data 0 0 32 0 INPUT NODEFVAL "data[31..0]"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @data 0 0 32 0 data 0 0 32 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL coshw.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL coshw.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL coshw.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL coshw.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL coshw_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
